module sigmo_lin32c(output signed [13:0] y, input signed [11:0] x);
wire [11:0] xabs = (x>=0) ? x : -x;
reg [14:0] f0, k;
always @* begin
    case (xabs[11:5])
    0: begin f0 = 8192; k = 16; end
    1: begin f0 = 8704; k = 16; end
    2: begin f0 = 9212; k = 16; end
    3: begin f0 = 9712; k = 15; end
    4: begin f0 = 10200; k = 15; end
    5: begin f0 = 10672; k = 14; end
    6: begin f0 = 11128; k = 14; end
    7: begin f0 = 11564; k = 13; end
    8: begin f0 = 11976; k = 12; end
    9: begin f0 = 12368; k = 12; end
    10: begin f0 = 12736; k = 11; end
    11: begin f0 = 13076; k = 10; end
    12: begin f0 = 13396; k = 9; end
    13: begin f0 = 13688; k = 8; end
    14: begin f0 = 13960; k = 8; end
    15: begin f0 = 14204; k = 7; end
    16: begin f0 = 14432; k = 6; end
    17: begin f0 = 14636; k = 6; end
    18: begin f0 = 14820; k = 5; end
    19: begin f0 = 14988; k = 5; end
    20: begin f0 = 15140; k = 4; end
    21: begin f0 = 15276; k = 4; end
    22: begin f0 = 15400; k = 3; end
    23: begin f0 = 15508; k = 3; end
    24: begin f0 = 15608; k = 3; end
    25: begin f0 = 15696; k = 2; end
    26: begin f0 = 15772; k = 2; end
    27: begin f0 = 15840; k = 2; end
    28: begin f0 = 15904; k = 2; end
    29: begin f0 = 15960; k = 2; end
    30: begin f0 = 16008; k = 1; end
    31: begin f0 = 16052; k = 1; end
    32: begin f0 = 16088; k = 1; end
    33: begin f0 = 16124; k = 1; end
    34: begin f0 = 16152; k = 1; end
    35: begin f0 = 16180; k = 1; end
    36: begin f0 = 16204; k = 1; end
    37: begin f0 = 16224; k = 1; end
    38: begin f0 = 16244; k = 0; end
    39: begin f0 = 16260; k = 0; end
    40: begin f0 = 16276; k = 0; end
    41: begin f0 = 16288; k = 0; end
    42: begin f0 = 16300; k = 0; end
    43: begin f0 = 16308; k = 0; end
    44: begin f0 = 16316; k = 0; end
    45: begin f0 = 16324; k = 0; end
    46: begin f0 = 16332; k = 0; end
    47: begin f0 = 16340; k = 0; end
    48: begin f0 = 16344; k = 0; end
    49: begin f0 = 16348; k = 0; end
    50: begin f0 = 16352; k = 0; end
    51: begin f0 = 16356; k = 0; end
    52: begin f0 = 16360; k = 0; end
    53: begin f0 = 16364; k = 0; end
    54: begin f0 = 16364; k = 0; end
    55: begin f0 = 16368; k = 0; end
    56: begin f0 = 16368; k = 0; end
    57: begin f0 = 16372; k = 0; end
    58: begin f0 = 16372; k = 0; end
    59: begin f0 = 16372; k = 0; end
    60: begin f0 = 16376; k = 0; end
    61: begin f0 = 16376; k = 0; end
    62: begin f0 = 16376; k = 0; end
    63: begin f0 = 16376; k = 0; end
    default: begin f0 = 16379; k = 0; end
    endcase
end
wire signed [15:0] yt0 = k*xabs[4:0] + f0;
wire signed [13:0] yt = yt0/4;
wire signed [3:0] diff;
compensation compensation (.diff(diff), .x(xabs[11:0]));
wire signed [13:0] yu = yt + {{10{diff[3]}},diff};
assign y = (x < 0) ? 4096 - yu : yu;
endmodule

module compensation (output reg signed [3:0] diff, input [11:0] x);
always @* begin
    case (x)
        0: diff =     0;
        1: diff =     0;
        2: diff =     0;
        3: diff =     0;
        4: diff =     0;
        5: diff =     0;
        6: diff =     0;
        7: diff =     0;
        8: diff =     0;
        9: diff =     0;
       10: diff =     0;
       11: diff =     0;
       12: diff =     0;
       13: diff =     0;
       14: diff =     0;
       15: diff =     0;
       16: diff =     0;
       17: diff =     0;
       18: diff =     0;
       19: diff =     0;
       20: diff =     0;
       21: diff =     0;
       22: diff =     0;
       23: diff =     0;
       24: diff =     0;
       25: diff =     0;
       26: diff =     0;
       27: diff =     0;
       28: diff =     0;
       29: diff =     0;
       30: diff =     0;
       31: diff =     0;
       32: diff =     0;
       33: diff =     0;
       34: diff =     0;
       35: diff =     0;
       36: diff =     0;
       37: diff =     0;
       38: diff =     0;
       39: diff =     0;
       40: diff =     0;
       41: diff =     0;
       42: diff =     0;
       43: diff =     0;
       44: diff =     0;
       45: diff =     0;
       46: diff =     0;
       47: diff =    -1;
       48: diff =    -1;
       49: diff =    -1;
       50: diff =    -1;
       51: diff =    -1;
       52: diff =    -1;
       53: diff =    -1;
       54: diff =    -1;
       55: diff =    -1;
       56: diff =    -1;
       57: diff =    -1;
       58: diff =    -1;
       59: diff =    -1;
       60: diff =    -1;
       61: diff =    -1;
       62: diff =    -1;
       63: diff =    -1;
       64: diff =     0;
       65: diff =     0;
       66: diff =     0;
       67: diff =    -1;
       68: diff =    -1;
       69: diff =    -1;
       70: diff =    -1;
       71: diff =    -1;
       72: diff =    -1;
       73: diff =    -1;
       74: diff =    -1;
       75: diff =    -1;
       76: diff =    -1;
       77: diff =    -1;
       78: diff =    -1;
       79: diff =    -1;
       80: diff =    -2;
       81: diff =    -2;
       82: diff =    -2;
       83: diff =    -2;
       84: diff =    -2;
       85: diff =    -2;
       86: diff =    -2;
       87: diff =    -2;
       88: diff =    -2;
       89: diff =    -3;
       90: diff =    -3;
       91: diff =    -3;
       92: diff =    -3;
       93: diff =    -3;
       94: diff =    -3;
       95: diff =    -3;
       96: diff =     0;
       97: diff =     0;
       98: diff =     0;
       99: diff =     0;
      100: diff =     0;
      101: diff =     1;
      102: diff =     1;
      103: diff =     1;
      104: diff =     0;
      105: diff =     1;
      106: diff =     1;
      107: diff =     1;
      108: diff =     1;
      109: diff =     2;
      110: diff =     1;
      111: diff =     1;
      112: diff =     1;
      113: diff =     2;
      114: diff =     2;
      115: diff =     1;
      116: diff =     1;
      117: diff =     2;
      118: diff =     2;
      119: diff =     2;
      120: diff =     1;
      121: diff =     2;
      122: diff =     2;
      123: diff =     2;
      124: diff =     2;
      125: diff =     2;
      126: diff =     2;
      127: diff =     2;
      128: diff =     0;
      129: diff =     0;
      130: diff =     0;
      131: diff =     0;
      132: diff =     0;
      133: diff =     0;
      134: diff =     0;
      135: diff =     0;
      136: diff =     0;
      137: diff =     0;
      138: diff =     0;
      139: diff =     0;
      140: diff =    -1;
      141: diff =     0;
      142: diff =     0;
      143: diff =     0;
      144: diff =    -1;
      145: diff =     0;
      146: diff =     0;
      147: diff =    -1;
      148: diff =    -1;
      149: diff =     0;
      150: diff =    -1;
      151: diff =    -1;
      152: diff =    -1;
      153: diff =    -1;
      154: diff =    -1;
      155: diff =    -1;
      156: diff =    -2;
      157: diff =    -1;
      158: diff =    -1;
      159: diff =    -2;
      160: diff =     0;
      161: diff =     1;
      162: diff =     0;
      163: diff =     1;
      164: diff =     0;
      165: diff =     1;
      166: diff =     1;
      167: diff =     1;
      168: diff =     1;
      169: diff =     1;
      170: diff =     1;
      171: diff =     2;
      172: diff =     1;
      173: diff =     2;
      174: diff =     1;
      175: diff =     2;
      176: diff =     2;
      177: diff =     2;
      178: diff =     2;
      179: diff =     2;
      180: diff =     2;
      181: diff =     2;
      182: diff =     2;
      183: diff =     2;
      184: diff =     2;
      185: diff =     2;
      186: diff =     2;
      187: diff =     2;
      188: diff =     2;
      189: diff =     2;
      190: diff =     2;
      191: diff =     2;
      192: diff =     0;
      193: diff =     0;
      194: diff =     0;
      195: diff =     0;
      196: diff =     0;
      197: diff =     0;
      198: diff =     0;
      199: diff =     0;
      200: diff =     0;
      201: diff =     0;
      202: diff =     0;
      203: diff =     0;
      204: diff =    -1;
      205: diff =     0;
      206: diff =    -1;
      207: diff =     0;
      208: diff =    -1;
      209: diff =    -1;
      210: diff =    -1;
      211: diff =    -1;
      212: diff =    -1;
      213: diff =    -1;
      214: diff =    -2;
      215: diff =    -1;
      216: diff =    -2;
      217: diff =    -1;
      218: diff =    -2;
      219: diff =    -2;
      220: diff =    -2;
      221: diff =    -2;
      222: diff =    -3;
      223: diff =    -2;
      224: diff =     0;
      225: diff =     0;
      226: diff =     1;
      227: diff =     1;
      228: diff =     0;
      229: diff =     0;
      230: diff =     1;
      231: diff =     1;
      232: diff =     0;
      233: diff =     1;
      234: diff =     1;
      235: diff =     1;
      236: diff =     0;
      237: diff =     1;
      238: diff =     1;
      239: diff =     1;
      240: diff =     0;
      241: diff =     1;
      242: diff =     1;
      243: diff =     1;
      244: diff =     0;
      245: diff =     0;
      246: diff =     1;
      247: diff =     1;
      248: diff =     0;
      249: diff =     0;
      250: diff =     0;
      251: diff =     1;
      252: diff =     0;
      253: diff =     0;
      254: diff =     0;
      255: diff =     0;
      256: diff =     0;
      257: diff =     1;
      258: diff =     1;
      259: diff =     1;
      260: diff =     1;
      261: diff =     1;
      262: diff =     1;
      263: diff =     1;
      264: diff =     1;
      265: diff =     1;
      266: diff =     2;
      267: diff =     2;
      268: diff =     2;
      269: diff =     2;
      270: diff =     2;
      271: diff =     2;
      272: diff =     2;
      273: diff =     2;
      274: diff =     2;
      275: diff =     2;
      276: diff =     2;
      277: diff =     2;
      278: diff =     2;
      279: diff =     2;
      280: diff =     2;
      281: diff =     2;
      282: diff =     2;
      283: diff =     2;
      284: diff =     2;
      285: diff =     2;
      286: diff =     2;
      287: diff =     2;
      288: diff =     0;
      289: diff =     0;
      290: diff =     0;
      291: diff =     0;
      292: diff =     0;
      293: diff =     0;
      294: diff =     0;
      295: diff =     0;
      296: diff =     0;
      297: diff =     0;
      298: diff =    -1;
      299: diff =    -1;
      300: diff =    -1;
      301: diff =    -1;
      302: diff =    -1;
      303: diff =    -1;
      304: diff =    -1;
      305: diff =    -1;
      306: diff =    -2;
      307: diff =    -2;
      308: diff =    -2;
      309: diff =    -2;
      310: diff =    -2;
      311: diff =    -2;
      312: diff =    -3;
      313: diff =    -3;
      314: diff =    -3;
      315: diff =    -3;
      316: diff =    -3;
      317: diff =    -4;
      318: diff =    -4;
      319: diff =    -4;
      320: diff =     0;
      321: diff =     1;
      322: diff =     0;
      323: diff =     0;
      324: diff =     0;
      325: diff =     1;
      326: diff =     0;
      327: diff =     0;
      328: diff =     0;
      329: diff =     1;
      330: diff =     0;
      331: diff =     0;
      332: diff =     0;
      333: diff =     0;
      334: diff =     0;
      335: diff =     0;
      336: diff =    -1;
      337: diff =     0;
      338: diff =     0;
      339: diff =    -1;
      340: diff =    -1;
      341: diff =     0;
      342: diff =    -1;
      343: diff =    -1;
      344: diff =    -1;
      345: diff =    -1;
      346: diff =    -1;
      347: diff =    -2;
      348: diff =    -2;
      349: diff =    -1;
      350: diff =    -2;
      351: diff =    -2;
      352: diff =     0;
      353: diff =     1;
      354: diff =     1;
      355: diff =     1;
      356: diff =     1;
      357: diff =     1;
      358: diff =     1;
      359: diff =     1;
      360: diff =     1;
      361: diff =     1;
      362: diff =     1;
      363: diff =     1;
      364: diff =     1;
      365: diff =     1;
      366: diff =     1;
      367: diff =     1;
      368: diff =     1;
      369: diff =     1;
      370: diff =     1;
      371: diff =     1;
      372: diff =     1;
      373: diff =     1;
      374: diff =     1;
      375: diff =     1;
      376: diff =     1;
      377: diff =     1;
      378: diff =     0;
      379: diff =     1;
      380: diff =     0;
      381: diff =     1;
      382: diff =     0;
      383: diff =     0;
      384: diff =     0;
      385: diff =     0;
      386: diff =     1;
      387: diff =     1;
      388: diff =     0;
      389: diff =     1;
      390: diff =     1;
      391: diff =     1;
      392: diff =     1;
      393: diff =     1;
      394: diff =     1;
      395: diff =     2;
      396: diff =     1;
      397: diff =     1;
      398: diff =     2;
      399: diff =     2;
      400: diff =     1;
      401: diff =     2;
      402: diff =     2;
      403: diff =     2;
      404: diff =     1;
      405: diff =     2;
      406: diff =     2;
      407: diff =     2;
      408: diff =     1;
      409: diff =     2;
      410: diff =     2;
      411: diff =     2;
      412: diff =     1;
      413: diff =     2;
      414: diff =     2;
      415: diff =     2;
      416: diff =     0;
      417: diff =     0;
      418: diff =     1;
      419: diff =     1;
      420: diff =     1;
      421: diff =     1;
      422: diff =     1;
      423: diff =     1;
      424: diff =     2;
      425: diff =     2;
      426: diff =     2;
      427: diff =     2;
      428: diff =     2;
      429: diff =     2;
      430: diff =     2;
      431: diff =     2;
      432: diff =     3;
      433: diff =     3;
      434: diff =     3;
      435: diff =     3;
      436: diff =     3;
      437: diff =     3;
      438: diff =     3;
      439: diff =     3;
      440: diff =     3;
      441: diff =     3;
      442: diff =     3;
      443: diff =     3;
      444: diff =     3;
      445: diff =     4;
      446: diff =     4;
      447: diff =     4;
      448: diff =     0;
      449: diff =     0;
      450: diff =     0;
      451: diff =     0;
      452: diff =     0;
      453: diff =     0;
      454: diff =     0;
      455: diff =     0;
      456: diff =     0;
      457: diff =     0;
      458: diff =     0;
      459: diff =    -1;
      460: diff =    -1;
      461: diff =    -1;
      462: diff =    -1;
      463: diff =    -1;
      464: diff =    -1;
      465: diff =    -1;
      466: diff =    -1;
      467: diff =    -1;
      468: diff =    -1;
      469: diff =    -1;
      470: diff =    -1;
      471: diff =    -1;
      472: diff =    -2;
      473: diff =    -2;
      474: diff =    -2;
      475: diff =    -2;
      476: diff =    -2;
      477: diff =    -2;
      478: diff =    -2;
      479: diff =    -2;
      480: diff =     0;
      481: diff =     1;
      482: diff =     1;
      483: diff =     1;
      484: diff =     1;
      485: diff =     2;
      486: diff =     1;
      487: diff =     1;
      488: diff =     1;
      489: diff =     2;
      490: diff =     2;
      491: diff =     1;
      492: diff =     1;
      493: diff =     2;
      494: diff =     2;
      495: diff =     1;
      496: diff =     1;
      497: diff =     2;
      498: diff =     2;
      499: diff =     1;
      500: diff =     1;
      501: diff =     2;
      502: diff =     2;
      503: diff =     1;
      504: diff =     1;
      505: diff =     2;
      506: diff =     2;
      507: diff =     1;
      508: diff =     1;
      509: diff =     2;
      510: diff =     1;
      511: diff =     1;
      512: diff =     0;
      513: diff =     0;
      514: diff =     0;
      515: diff =     1;
      516: diff =     0;
      517: diff =     1;
      518: diff =     1;
      519: diff =     1;
      520: diff =     1;
      521: diff =     2;
      522: diff =     1;
      523: diff =     2;
      524: diff =     2;
      525: diff =     2;
      526: diff =     2;
      527: diff =     2;
      528: diff =     2;
      529: diff =     3;
      530: diff =     2;
      531: diff =     3;
      532: diff =     2;
      533: diff =     3;
      534: diff =     3;
      535: diff =     3;
      536: diff =     3;
      537: diff =     3;
      538: diff =     3;
      539: diff =     3;
      540: diff =     3;
      541: diff =     3;
      542: diff =     3;
      543: diff =     3;
      544: diff =     0;
      545: diff =     1;
      546: diff =     0;
      547: diff =     1;
      548: diff =     0;
      549: diff =     1;
      550: diff =     0;
      551: diff =     1;
      552: diff =     0;
      553: diff =     1;
      554: diff =     0;
      555: diff =     0;
      556: diff =     0;
      557: diff =     0;
      558: diff =     0;
      559: diff =     0;
      560: diff =     0;
      561: diff =     0;
      562: diff =     0;
      563: diff =     0;
      564: diff =     0;
      565: diff =     0;
      566: diff =    -1;
      567: diff =     0;
      568: diff =    -1;
      569: diff =     0;
      570: diff =    -1;
      571: diff =    -1;
      572: diff =    -1;
      573: diff =    -1;
      574: diff =    -1;
      575: diff =    -1;
      576: diff =     0;
      577: diff =     1;
      578: diff =     1;
      579: diff =     2;
      580: diff =     1;
      581: diff =     1;
      582: diff =     2;
      583: diff =     2;
      584: diff =     1;
      585: diff =     2;
      586: diff =     2;
      587: diff =     2;
      588: diff =     2;
      589: diff =     2;
      590: diff =     2;
      591: diff =     3;
      592: diff =     2;
      593: diff =     2;
      594: diff =     3;
      595: diff =     3;
      596: diff =     2;
      597: diff =     2;
      598: diff =     3;
      599: diff =     3;
      600: diff =     2;
      601: diff =     3;
      602: diff =     3;
      603: diff =     3;
      604: diff =     2;
      605: diff =     3;
      606: diff =     3;
      607: diff =     3;
      608: diff =     0;
      609: diff =     1;
      610: diff =     1;
      611: diff =     1;
      612: diff =     0;
      613: diff =     1;
      614: diff =     1;
      615: diff =     1;
      616: diff =     0;
      617: diff =     0;
      618: diff =     1;
      619: diff =     1;
      620: diff =     0;
      621: diff =     0;
      622: diff =     0;
      623: diff =     1;
      624: diff =     0;
      625: diff =     0;
      626: diff =     0;
      627: diff =     0;
      628: diff =     0;
      629: diff =     0;
      630: diff =     0;
      631: diff =     0;
      632: diff =    -1;
      633: diff =    -1;
      634: diff =    -1;
      635: diff =     0;
      636: diff =    -1;
      637: diff =    -1;
      638: diff =    -1;
      639: diff =    -1;
      640: diff =     0;
      641: diff =     0;
      642: diff =     1;
      643: diff =     1;
      644: diff =     1;
      645: diff =     1;
      646: diff =     1;
      647: diff =     1;
      648: diff =     1;
      649: diff =     1;
      650: diff =     1;
      651: diff =     1;
      652: diff =     1;
      653: diff =     2;
      654: diff =     2;
      655: diff =     2;
      656: diff =     2;
      657: diff =     2;
      658: diff =     2;
      659: diff =     2;
      660: diff =     2;
      661: diff =     2;
      662: diff =     2;
      663: diff =     2;
      664: diff =     2;
      665: diff =     2;
      666: diff =     2;
      667: diff =     2;
      668: diff =     2;
      669: diff =     2;
      670: diff =     2;
      671: diff =     2;
      672: diff =     0;
      673: diff =     0;
      674: diff =     0;
      675: diff =     0;
      676: diff =     0;
      677: diff =     0;
      678: diff =     0;
      679: diff =     0;
      680: diff =     0;
      681: diff =     0;
      682: diff =     0;
      683: diff =     0;
      684: diff =     0;
      685: diff =     0;
      686: diff =     0;
      687: diff =     0;
      688: diff =     0;
      689: diff =     0;
      690: diff =     0;
      691: diff =     0;
      692: diff =     0;
      693: diff =     0;
      694: diff =     0;
      695: diff =     0;
      696: diff =     0;
      697: diff =    -1;
      698: diff =    -1;
      699: diff =    -1;
      700: diff =    -1;
      701: diff =    -1;
      702: diff =    -1;
      703: diff =    -1;
      704: diff =     0;
      705: diff =     1;
      706: diff =     1;
      707: diff =     1;
      708: diff =     0;
      709: diff =     1;
      710: diff =     1;
      711: diff =     1;
      712: diff =     1;
      713: diff =     2;
      714: diff =     2;
      715: diff =     2;
      716: diff =     2;
      717: diff =     2;
      718: diff =     2;
      719: diff =     2;
      720: diff =     2;
      721: diff =     3;
      722: diff =     3;
      723: diff =     3;
      724: diff =     2;
      725: diff =     3;
      726: diff =     3;
      727: diff =     3;
      728: diff =     3;
      729: diff =     4;
      730: diff =     3;
      731: diff =     3;
      732: diff =     3;
      733: diff =     4;
      734: diff =     4;
      735: diff =     3;
      736: diff =     0;
      737: diff =     1;
      738: diff =     1;
      739: diff =     1;
      740: diff =     0;
      741: diff =     1;
      742: diff =     1;
      743: diff =     1;
      744: diff =     1;
      745: diff =     1;
      746: diff =     1;
      747: diff =     1;
      748: diff =     1;
      749: diff =     2;
      750: diff =     1;
      751: diff =     1;
      752: diff =     1;
      753: diff =     2;
      754: diff =     1;
      755: diff =     1;
      756: diff =     1;
      757: diff =     2;
      758: diff =     1;
      759: diff =     1;
      760: diff =     1;
      761: diff =     2;
      762: diff =     1;
      763: diff =     1;
      764: diff =     1;
      765: diff =     2;
      766: diff =     1;
      767: diff =     1;
      768: diff =     0;
      769: diff =     0;
      770: diff =     0;
      771: diff =     0;
      772: diff =     0;
      773: diff =     0;
      774: diff =     0;
      775: diff =     0;
      776: diff =    -1;
      777: diff =     0;
      778: diff =     0;
      779: diff =     0;
      780: diff =    -1;
      781: diff =     0;
      782: diff =     0;
      783: diff =    -1;
      784: diff =    -1;
      785: diff =     0;
      786: diff =    -1;
      787: diff =    -1;
      788: diff =    -1;
      789: diff =    -1;
      790: diff =    -1;
      791: diff =    -1;
      792: diff =    -2;
      793: diff =    -1;
      794: diff =    -1;
      795: diff =    -2;
      796: diff =    -2;
      797: diff =    -1;
      798: diff =    -2;
      799: diff =    -2;
      800: diff =     0;
      801: diff =     0;
      802: diff =     0;
      803: diff =     1;
      804: diff =     0;
      805: diff =     1;
      806: diff =     0;
      807: diff =     1;
      808: diff =     1;
      809: diff =     1;
      810: diff =     1;
      811: diff =     2;
      812: diff =     1;
      813: diff =     2;
      814: diff =     1;
      815: diff =     2;
      816: diff =     2;
      817: diff =     2;
      818: diff =     2;
      819: diff =     2;
      820: diff =     2;
      821: diff =     3;
      822: diff =     2;
      823: diff =     3;
      824: diff =     2;
      825: diff =     3;
      826: diff =     3;
      827: diff =     3;
      828: diff =     3;
      829: diff =     3;
      830: diff =     3;
      831: diff =     4;
      832: diff =     0;
      833: diff =     1;
      834: diff =     0;
      835: diff =     1;
      836: diff =     0;
      837: diff =     1;
      838: diff =     1;
      839: diff =     1;
      840: diff =     1;
      841: diff =     1;
      842: diff =     1;
      843: diff =     1;
      844: diff =     1;
      845: diff =     1;
      846: diff =     1;
      847: diff =     2;
      848: diff =     1;
      849: diff =     2;
      850: diff =     1;
      851: diff =     2;
      852: diff =     1;
      853: diff =     2;
      854: diff =     1;
      855: diff =     2;
      856: diff =     1;
      857: diff =     2;
      858: diff =     1;
      859: diff =     2;
      860: diff =     1;
      861: diff =     2;
      862: diff =     1;
      863: diff =     2;
      864: diff =     0;
      865: diff =     1;
      866: diff =     0;
      867: diff =     1;
      868: diff =     1;
      869: diff =     1;
      870: diff =     1;
      871: diff =     1;
      872: diff =     1;
      873: diff =     1;
      874: diff =     1;
      875: diff =     1;
      876: diff =     0;
      877: diff =     1;
      878: diff =     0;
      879: diff =     1;
      880: diff =     0;
      881: diff =     1;
      882: diff =     0;
      883: diff =     1;
      884: diff =     0;
      885: diff =     1;
      886: diff =     0;
      887: diff =     1;
      888: diff =     0;
      889: diff =     1;
      890: diff =     0;
      891: diff =     1;
      892: diff =     0;
      893: diff =     1;
      894: diff =     0;
      895: diff =     0;
      896: diff =     0;
      897: diff =     0;
      898: diff =     0;
      899: diff =     0;
      900: diff =     0;
      901: diff =     0;
      902: diff =     0;
      903: diff =     0;
      904: diff =     0;
      905: diff =     0;
      906: diff =    -1;
      907: diff =     0;
      908: diff =    -1;
      909: diff =     0;
      910: diff =    -1;
      911: diff =     0;
      912: diff =    -1;
      913: diff =    -1;
      914: diff =    -1;
      915: diff =    -1;
      916: diff =    -1;
      917: diff =    -1;
      918: diff =    -1;
      919: diff =    -1;
      920: diff =    -2;
      921: diff =    -1;
      922: diff =    -2;
      923: diff =    -1;
      924: diff =    -2;
      925: diff =    -2;
      926: diff =    -2;
      927: diff =    -2;
      928: diff =     0;
      929: diff =     0;
      930: diff =    -1;
      931: diff =     0;
      932: diff =    -1;
      933: diff =     0;
      934: diff =    -1;
      935: diff =    -1;
      936: diff =    -1;
      937: diff =    -1;
      938: diff =    -1;
      939: diff =    -1;
      940: diff =    -2;
      941: diff =    -1;
      942: diff =    -2;
      943: diff =    -1;
      944: diff =    -2;
      945: diff =    -2;
      946: diff =    -2;
      947: diff =    -2;
      948: diff =    -3;
      949: diff =    -2;
      950: diff =    -3;
      951: diff =    -2;
      952: diff =    -3;
      953: diff =    -3;
      954: diff =    -3;
      955: diff =    -3;
      956: diff =    -4;
      957: diff =    -3;
      958: diff =    -4;
      959: diff =    -3;
      960: diff =     0;
      961: diff =     0;
      962: diff =     1;
      963: diff =     1;
      964: diff =     0;
      965: diff =     1;
      966: diff =     1;
      967: diff =     1;
      968: diff =     1;
      969: diff =     1;
      970: diff =     1;
      971: diff =     2;
      972: diff =     1;
      973: diff =     1;
      974: diff =     2;
      975: diff =     2;
      976: diff =     1;
      977: diff =     2;
      978: diff =     2;
      979: diff =     2;
      980: diff =     2;
      981: diff =     2;
      982: diff =     2;
      983: diff =     3;
      984: diff =     2;
      985: diff =     2;
      986: diff =     3;
      987: diff =     3;
      988: diff =     2;
      989: diff =     3;
      990: diff =     3;
      991: diff =     3;
      992: diff =     0;
      993: diff =     0;
      994: diff =     0;
      995: diff =     1;
      996: diff =     0;
      997: diff =     0;
      998: diff =     1;
      999: diff =     1;
     1000: diff =     0;
     1001: diff =     1;
     1002: diff =     1;
     1003: diff =     1;
     1004: diff =     0;
     1005: diff =     1;
     1006: diff =     1;
     1007: diff =     1;
     1008: diff =     1;
     1009: diff =     1;
     1010: diff =     1;
     1011: diff =     2;
     1012: diff =     1;
     1013: diff =     1;
     1014: diff =     1;
     1015: diff =     2;
     1016: diff =     1;
     1017: diff =     1;
     1018: diff =     2;
     1019: diff =     2;
     1020: diff =     1;
     1021: diff =     1;
     1022: diff =     2;
     1023: diff =     2;
     1024: diff =     0;
     1025: diff =     1;
     1026: diff =     1;
     1027: diff =     1;
     1028: diff =     0;
     1029: diff =     1;
     1030: diff =     1;
     1031: diff =     1;
     1032: diff =     1;
     1033: diff =     1;
     1034: diff =     1;
     1035: diff =     1;
     1036: diff =     1;
     1037: diff =     1;
     1038: diff =     1;
     1039: diff =     1;
     1040: diff =     1;
     1041: diff =     1;
     1042: diff =     1;
     1043: diff =     2;
     1044: diff =     1;
     1045: diff =     1;
     1046: diff =     1;
     1047: diff =     2;
     1048: diff =     1;
     1049: diff =     1;
     1050: diff =     1;
     1051: diff =     2;
     1052: diff =     1;
     1053: diff =     1;
     1054: diff =     1;
     1055: diff =     2;
     1056: diff =     0;
     1057: diff =     0;
     1058: diff =     0;
     1059: diff =     1;
     1060: diff =     0;
     1061: diff =     0;
     1062: diff =     0;
     1063: diff =     1;
     1064: diff =     0;
     1065: diff =     0;
     1066: diff =     0;
     1067: diff =     1;
     1068: diff =     0;
     1069: diff =     0;
     1070: diff =     0;
     1071: diff =     0;
     1072: diff =     0;
     1073: diff =     0;
     1074: diff =     0;
     1075: diff =     0;
     1076: diff =     0;
     1077: diff =     0;
     1078: diff =     0;
     1079: diff =     0;
     1080: diff =     0;
     1081: diff =     0;
     1082: diff =     0;
     1083: diff =     0;
     1084: diff =     0;
     1085: diff =     0;
     1086: diff =     0;
     1087: diff =     0;
     1088: diff =     0;
     1089: diff =     1;
     1090: diff =     1;
     1091: diff =     1;
     1092: diff =     0;
     1093: diff =     0;
     1094: diff =     1;
     1095: diff =     1;
     1096: diff =     0;
     1097: diff =     0;
     1098: diff =     1;
     1099: diff =     1;
     1100: diff =     0;
     1101: diff =     0;
     1102: diff =     0;
     1103: diff =     1;
     1104: diff =     0;
     1105: diff =     0;
     1106: diff =     0;
     1107: diff =     0;
     1108: diff =     0;
     1109: diff =     0;
     1110: diff =     0;
     1111: diff =     0;
     1112: diff =    -1;
     1113: diff =     0;
     1114: diff =     0;
     1115: diff =     0;
     1116: diff =    -1;
     1117: diff =    -1;
     1118: diff =     0;
     1119: diff =     0;
     1120: diff =     0;
     1121: diff =     0;
     1122: diff =     0;
     1123: diff =     1;
     1124: diff =     0;
     1125: diff =     0;
     1126: diff =     0;
     1127: diff =     0;
     1128: diff =     0;
     1129: diff =     0;
     1130: diff =     0;
     1131: diff =     0;
     1132: diff =    -1;
     1133: diff =     0;
     1134: diff =     0;
     1135: diff =     0;
     1136: diff =    -1;
     1137: diff =    -1;
     1138: diff =    -1;
     1139: diff =     0;
     1140: diff =    -1;
     1141: diff =    -1;
     1142: diff =    -1;
     1143: diff =    -1;
     1144: diff =    -1;
     1145: diff =    -1;
     1146: diff =    -1;
     1147: diff =    -1;
     1148: diff =    -2;
     1149: diff =    -2;
     1150: diff =    -1;
     1151: diff =    -1;
     1152: diff =     0;
     1153: diff =     0;
     1154: diff =     0;
     1155: diff =     1;
     1156: diff =     0;
     1157: diff =     0;
     1158: diff =     0;
     1159: diff =     0;
     1160: diff =    -1;
     1161: diff =     0;
     1162: diff =     0;
     1163: diff =     0;
     1164: diff =    -1;
     1165: diff =    -1;
     1166: diff =    -1;
     1167: diff =     0;
     1168: diff =    -1;
     1169: diff =    -1;
     1170: diff =    -1;
     1171: diff =    -1;
     1172: diff =    -2;
     1173: diff =    -1;
     1174: diff =    -1;
     1175: diff =    -1;
     1176: diff =    -2;
     1177: diff =    -2;
     1178: diff =    -2;
     1179: diff =    -2;
     1180: diff =    -2;
     1181: diff =    -2;
     1182: diff =    -2;
     1183: diff =    -2;
     1184: diff =     0;
     1185: diff =     0;
     1186: diff =     1;
     1187: diff =     1;
     1188: diff =     0;
     1189: diff =     0;
     1190: diff =     0;
     1191: diff =     0;
     1192: diff =    -1;
     1193: diff =     0;
     1194: diff =     0;
     1195: diff =     0;
     1196: diff =    -1;
     1197: diff =    -1;
     1198: diff =    -1;
     1199: diff =    -1;
     1200: diff =    -1;
     1201: diff =    -1;
     1202: diff =    -1;
     1203: diff =    -1;
     1204: diff =    -2;
     1205: diff =    -2;
     1206: diff =    -2;
     1207: diff =    -1;
     1208: diff =    -2;
     1209: diff =    -2;
     1210: diff =    -2;
     1211: diff =    -2;
     1212: diff =    -3;
     1213: diff =    -3;
     1214: diff =    -2;
     1215: diff =    -2;
     1216: diff =     0;
     1217: diff =     0;
     1218: diff =     0;
     1219: diff =     0;
     1220: diff =     0;
     1221: diff =     1;
     1222: diff =     1;
     1223: diff =     1;
     1224: diff =     1;
     1225: diff =     1;
     1226: diff =     1;
     1227: diff =     1;
     1228: diff =     1;
     1229: diff =     2;
     1230: diff =     2;
     1231: diff =     2;
     1232: diff =     2;
     1233: diff =     2;
     1234: diff =     2;
     1235: diff =     2;
     1236: diff =     2;
     1237: diff =     3;
     1238: diff =     3;
     1239: diff =     3;
     1240: diff =     3;
     1241: diff =     3;
     1242: diff =     3;
     1243: diff =     3;
     1244: diff =     3;
     1245: diff =     4;
     1246: diff =     4;
     1247: diff =     4;
     1248: diff =     0;
     1249: diff =     0;
     1250: diff =     0;
     1251: diff =     0;
     1252: diff =     0;
     1253: diff =     1;
     1254: diff =     1;
     1255: diff =     1;
     1256: diff =     1;
     1257: diff =     1;
     1258: diff =     1;
     1259: diff =     1;
     1260: diff =     1;
     1261: diff =     1;
     1262: diff =     2;
     1263: diff =     2;
     1264: diff =     2;
     1265: diff =     2;
     1266: diff =     2;
     1267: diff =     2;
     1268: diff =     2;
     1269: diff =     2;
     1270: diff =     3;
     1271: diff =     3;
     1272: diff =     3;
     1273: diff =     3;
     1274: diff =     3;
     1275: diff =     3;
     1276: diff =     3;
     1277: diff =     3;
     1278: diff =     3;
     1279: diff =     3;
     1280: diff =     0;
     1281: diff =     0;
     1282: diff =     0;
     1283: diff =     0;
     1284: diff =     0;
     1285: diff =     0;
     1286: diff =     0;
     1287: diff =     0;
     1288: diff =     0;
     1289: diff =     1;
     1290: diff =     1;
     1291: diff =     1;
     1292: diff =     1;
     1293: diff =     1;
     1294: diff =     1;
     1295: diff =     1;
     1296: diff =     1;
     1297: diff =     1;
     1298: diff =     1;
     1299: diff =     2;
     1300: diff =     2;
     1301: diff =     2;
     1302: diff =     2;
     1303: diff =     2;
     1304: diff =     2;
     1305: diff =     2;
     1306: diff =     2;
     1307: diff =     2;
     1308: diff =     2;
     1309: diff =     3;
     1310: diff =     3;
     1311: diff =     3;
     1312: diff =     0;
     1313: diff =     0;
     1314: diff =     0;
     1315: diff =     0;
     1316: diff =     0;
     1317: diff =     0;
     1318: diff =     0;
     1319: diff =     0;
     1320: diff =     1;
     1321: diff =     1;
     1322: diff =     1;
     1323: diff =     1;
     1324: diff =     1;
     1325: diff =     1;
     1326: diff =     1;
     1327: diff =     1;
     1328: diff =     1;
     1329: diff =     1;
     1330: diff =     1;
     1331: diff =     2;
     1332: diff =     2;
     1333: diff =     2;
     1334: diff =     2;
     1335: diff =     2;
     1336: diff =     2;
     1337: diff =     2;
     1338: diff =     2;
     1339: diff =     2;
     1340: diff =     2;
     1341: diff =     2;
     1342: diff =     2;
     1343: diff =     3;
     1344: diff =     0;
     1345: diff =     0;
     1346: diff =     0;
     1347: diff =     0;
     1348: diff =     0;
     1349: diff =     0;
     1350: diff =     0;
     1351: diff =     0;
     1352: diff =     0;
     1353: diff =     0;
     1354: diff =     0;
     1355: diff =     1;
     1356: diff =     1;
     1357: diff =     1;
     1358: diff =     1;
     1359: diff =     1;
     1360: diff =     1;
     1361: diff =     1;
     1362: diff =     1;
     1363: diff =     1;
     1364: diff =     1;
     1365: diff =     1;
     1366: diff =     1;
     1367: diff =     1;
     1368: diff =     2;
     1369: diff =     2;
     1370: diff =     2;
     1371: diff =     2;
     1372: diff =     2;
     1373: diff =     2;
     1374: diff =     2;
     1375: diff =     2;
     1376: diff =     0;
     1377: diff =     0;
     1378: diff =     0;
     1379: diff =     0;
     1380: diff =     0;
     1381: diff =     0;
     1382: diff =     1;
     1383: diff =     1;
     1384: diff =     1;
     1385: diff =     1;
     1386: diff =     1;
     1387: diff =     1;
     1388: diff =     1;
     1389: diff =     1;
     1390: diff =     1;
     1391: diff =     1;
     1392: diff =     1;
     1393: diff =     1;
     1394: diff =     1;
     1395: diff =     1;
     1396: diff =     2;
     1397: diff =     2;
     1398: diff =     2;
     1399: diff =     2;
     1400: diff =     2;
     1401: diff =     2;
     1402: diff =     2;
     1403: diff =     2;
     1404: diff =     2;
     1405: diff =     2;
     1406: diff =     2;
     1407: diff =     2;
     1408: diff =     0;
     1409: diff =     0;
     1410: diff =     0;
     1411: diff =     1;
     1412: diff =     1;
     1413: diff =     1;
     1414: diff =     1;
     1415: diff =     1;
     1416: diff =     1;
     1417: diff =     1;
     1418: diff =     1;
     1419: diff =     1;
     1420: diff =     1;
     1421: diff =     1;
     1422: diff =     1;
     1423: diff =     1;
     1424: diff =     1;
     1425: diff =     1;
     1426: diff =     1;
     1427: diff =     2;
     1428: diff =     2;
     1429: diff =     2;
     1430: diff =     2;
     1431: diff =     2;
     1432: diff =     2;
     1433: diff =     2;
     1434: diff =     2;
     1435: diff =     2;
     1436: diff =     2;
     1437: diff =     2;
     1438: diff =     2;
     1439: diff =     2;
     1440: diff =     0;
     1441: diff =     0;
     1442: diff =     0;
     1443: diff =     0;
     1444: diff =     1;
     1445: diff =     1;
     1446: diff =     1;
     1447: diff =     1;
     1448: diff =     1;
     1449: diff =     1;
     1450: diff =     1;
     1451: diff =     1;
     1452: diff =     1;
     1453: diff =     1;
     1454: diff =     1;
     1455: diff =     1;
     1456: diff =     1;
     1457: diff =     1;
     1458: diff =     1;
     1459: diff =     1;
     1460: diff =     1;
     1461: diff =     1;
     1462: diff =     1;
     1463: diff =     2;
     1464: diff =     2;
     1465: diff =     2;
     1466: diff =     2;
     1467: diff =     2;
     1468: diff =     2;
     1469: diff =     2;
     1470: diff =     2;
     1471: diff =     2;
     1472: diff =     0;
     1473: diff =     0;
     1474: diff =     0;
     1475: diff =     0;
     1476: diff =     0;
     1477: diff =     0;
     1478: diff =     0;
     1479: diff =     0;
     1480: diff =     0;
     1481: diff =     0;
     1482: diff =     1;
     1483: diff =     1;
     1484: diff =     1;
     1485: diff =     1;
     1486: diff =     1;
     1487: diff =     1;
     1488: diff =     1;
     1489: diff =     1;
     1490: diff =     1;
     1491: diff =     1;
     1492: diff =     1;
     1493: diff =     1;
     1494: diff =     1;
     1495: diff =     1;
     1496: diff =     1;
     1497: diff =     1;
     1498: diff =     1;
     1499: diff =     1;
     1500: diff =     1;
     1501: diff =     1;
     1502: diff =     1;
     1503: diff =     1;
     1504: diff =     0;
     1505: diff =     0;
     1506: diff =     0;
     1507: diff =     0;
     1508: diff =     0;
     1509: diff =     0;
     1510: diff =     0;
     1511: diff =     0;
     1512: diff =     0;
     1513: diff =     0;
     1514: diff =     0;
     1515: diff =     0;
     1516: diff =     0;
     1517: diff =     0;
     1518: diff =     0;
     1519: diff =     0;
     1520: diff =     0;
     1521: diff =     0;
     1522: diff =     0;
     1523: diff =     0;
     1524: diff =     0;
     1525: diff =     0;
     1526: diff =     0;
     1527: diff =     1;
     1528: diff =     1;
     1529: diff =     1;
     1530: diff =     1;
     1531: diff =     1;
     1532: diff =     1;
     1533: diff =     1;
     1534: diff =     1;
     1535: diff =     1;
     1536: diff =     0;
     1537: diff =     0;
     1538: diff =     0;
     1539: diff =     0;
     1540: diff =     0;
     1541: diff =     0;
     1542: diff =     0;
     1543: diff =     0;
     1544: diff =     0;
     1545: diff =     0;
     1546: diff =     0;
     1547: diff =     0;
     1548: diff =     0;
     1549: diff =     0;
     1550: diff =     0;
     1551: diff =     0;
     1552: diff =     0;
     1553: diff =     1;
     1554: diff =     1;
     1555: diff =     1;
     1556: diff =     1;
     1557: diff =     1;
     1558: diff =     1;
     1559: diff =     1;
     1560: diff =     1;
     1561: diff =     1;
     1562: diff =     1;
     1563: diff =     1;
     1564: diff =     1;
     1565: diff =     1;
     1566: diff =     1;
     1567: diff =     1;
     1568: diff =     0;
     1569: diff =     0;
     1570: diff =     0;
     1571: diff =     0;
     1572: diff =     0;
     1573: diff =     0;
     1574: diff =     0;
     1575: diff =     0;
     1576: diff =     0;
     1577: diff =     0;
     1578: diff =     0;
     1579: diff =     0;
     1580: diff =     0;
     1581: diff =     1;
     1582: diff =     1;
     1583: diff =     1;
     1584: diff =     1;
     1585: diff =     1;
     1586: diff =     1;
     1587: diff =     1;
     1588: diff =     1;
     1589: diff =     1;
     1590: diff =     1;
     1591: diff =     1;
     1592: diff =     1;
     1593: diff =     1;
     1594: diff =     1;
     1595: diff =     1;
     1596: diff =     1;
     1597: diff =     1;
     1598: diff =     1;
     1599: diff =     1;
     1600: diff =     0;
     1601: diff =     0;
     1602: diff =     0;
     1603: diff =     0;
     1604: diff =     0;
     1605: diff =     0;
     1606: diff =     0;
     1607: diff =     0;
     1608: diff =     0;
     1609: diff =     0;
     1610: diff =     0;
     1611: diff =     0;
     1612: diff =     0;
     1613: diff =     0;
     1614: diff =     1;
     1615: diff =     1;
     1616: diff =     1;
     1617: diff =     1;
     1618: diff =     1;
     1619: diff =     1;
     1620: diff =     1;
     1621: diff =     1;
     1622: diff =     1;
     1623: diff =     1;
     1624: diff =     1;
     1625: diff =     1;
     1626: diff =     1;
     1627: diff =     1;
     1628: diff =     1;
     1629: diff =     1;
     1630: diff =     1;
     1631: diff =     1;
     1632: diff =     0;
     1633: diff =     0;
     1634: diff =     0;
     1635: diff =     0;
     1636: diff =     0;
     1637: diff =     0;
     1638: diff =     0;
     1639: diff =     0;
     1640: diff =     0;
     1641: diff =     0;
     1642: diff =     0;
     1643: diff =     0;
     1644: diff =     0;
     1645: diff =     0;
     1646: diff =     0;
     1647: diff =     0;
     1648: diff =     0;
     1649: diff =     0;
     1650: diff =     1;
     1651: diff =     1;
     1652: diff =     1;
     1653: diff =     1;
     1654: diff =     1;
     1655: diff =     1;
     1656: diff =     1;
     1657: diff =     1;
     1658: diff =     1;
     1659: diff =     1;
     1660: diff =     1;
     1661: diff =     1;
     1662: diff =     1;
     1663: diff =     1;
     1664: diff =     0;
     1665: diff =     0;
     1666: diff =     0;
     1667: diff =     0;
     1668: diff =     0;
     1669: diff =     0;
     1670: diff =     0;
     1671: diff =     0;
     1672: diff =     0;
     1673: diff =     0;
     1674: diff =     0;
     1675: diff =     0;
     1676: diff =     0;
     1677: diff =     0;
     1678: diff =     0;
     1679: diff =     0;
     1680: diff =     0;
     1681: diff =     0;
     1682: diff =     0;
     1683: diff =     0;
     1684: diff =     0;
     1685: diff =     0;
     1686: diff =     0;
     1687: diff =     0;
     1688: diff =     0;
     1689: diff =     0;
     1690: diff =     0;
     1691: diff =     0;
     1692: diff =     0;
     1693: diff =     1;
     1694: diff =     1;
     1695: diff =     1;
     1696: diff =     0;
     1697: diff =     0;
     1698: diff =     0;
     1699: diff =     0;
     1700: diff =     0;
     1701: diff =     0;
     1702: diff =     0;
     1703: diff =     0;
     1704: diff =     0;
     1705: diff =     0;
     1706: diff =     0;
     1707: diff =     0;
     1708: diff =     0;
     1709: diff =     0;
     1710: diff =     0;
     1711: diff =     0;
     1712: diff =     0;
     1713: diff =     0;
     1714: diff =     0;
     1715: diff =     0;
     1716: diff =     0;
     1717: diff =     0;
     1718: diff =     0;
     1719: diff =     0;
     1720: diff =     0;
     1721: diff =     0;
     1722: diff =     0;
     1723: diff =     0;
     1724: diff =     0;
     1725: diff =     0;
     1726: diff =     0;
     1727: diff =     0;
     1728: diff =     0;
     1729: diff =     0;
     1730: diff =     0;
     1731: diff =     0;
     1732: diff =     0;
     1733: diff =     0;
     1734: diff =     0;
     1735: diff =     0;
     1736: diff =     0;
     1737: diff =     0;
     1738: diff =     0;
     1739: diff =     0;
     1740: diff =     0;
     1741: diff =     0;
     1742: diff =     0;
     1743: diff =     0;
     1744: diff =     0;
     1745: diff =     1;
     1746: diff =     1;
     1747: diff =     1;
     1748: diff =     1;
     1749: diff =     1;
     1750: diff =     1;
     1751: diff =     1;
     1752: diff =     1;
     1753: diff =     1;
     1754: diff =     1;
     1755: diff =     1;
     1756: diff =     1;
     1757: diff =     1;
     1758: diff =     1;
     1759: diff =     1;
     1760: diff =     0;
     1761: diff =     0;
     1762: diff =     0;
     1763: diff =     0;
     1764: diff =     0;
     1765: diff =     0;
     1766: diff =     0;
     1767: diff =     0;
     1768: diff =     0;
     1769: diff =     0;
     1770: diff =     0;
     1771: diff =     0;
     1772: diff =     0;
     1773: diff =     0;
     1774: diff =     0;
     1775: diff =     0;
     1776: diff =     0;
     1777: diff =     0;
     1778: diff =     0;
     1779: diff =     0;
     1780: diff =     0;
     1781: diff =     0;
     1782: diff =     0;
     1783: diff =     0;
     1784: diff =     0;
     1785: diff =     0;
     1786: diff =     0;
     1787: diff =     0;
     1788: diff =     0;
     1789: diff =     0;
     1790: diff =     0;
     1791: diff =     0;
     1792: diff =     0;
     1793: diff =     0;
     1794: diff =     0;
     1795: diff =     0;
     1796: diff =     0;
     1797: diff =     0;
     1798: diff =     0;
     1799: diff =     0;
     1800: diff =     0;
     1801: diff =     0;
     1802: diff =     0;
     1803: diff =     0;
     1804: diff =     0;
     1805: diff =     0;
     1806: diff =     0;
     1807: diff =     0;
     1808: diff =     0;
     1809: diff =     1;
     1810: diff =     1;
     1811: diff =     1;
     1812: diff =     1;
     1813: diff =     1;
     1814: diff =     1;
     1815: diff =     1;
     1816: diff =     1;
     1817: diff =     1;
     1818: diff =     1;
     1819: diff =     1;
     1820: diff =     1;
     1821: diff =     1;
     1822: diff =     1;
     1823: diff =     1;
     1824: diff =     0;
     1825: diff =     0;
     1826: diff =     0;
     1827: diff =     0;
     1828: diff =     0;
     1829: diff =     0;
     1830: diff =     0;
     1831: diff =     0;
     1832: diff =     0;
     1833: diff =     0;
     1834: diff =     0;
     1835: diff =     0;
     1836: diff =     0;
     1837: diff =     0;
     1838: diff =     0;
     1839: diff =     0;
     1840: diff =     0;
     1841: diff =     0;
     1842: diff =     0;
     1843: diff =     0;
     1844: diff =     0;
     1845: diff =     0;
     1846: diff =     0;
     1847: diff =     0;
     1848: diff =     0;
     1849: diff =     0;
     1850: diff =     0;
     1851: diff =     0;
     1852: diff =     0;
     1853: diff =     0;
     1854: diff =     0;
     1855: diff =     0;
     1856: diff =     0;
     1857: diff =     0;
     1858: diff =     0;
     1859: diff =     0;
     1860: diff =     0;
     1861: diff =     0;
     1862: diff =     0;
     1863: diff =     0;
     1864: diff =     0;
     1865: diff =     0;
     1866: diff =     0;
     1867: diff =     0;
     1868: diff =     0;
     1869: diff =     0;
     1870: diff =     0;
     1871: diff =     0;
     1872: diff =     0;
     1873: diff =     0;
     1874: diff =     0;
     1875: diff =     0;
     1876: diff =     0;
     1877: diff =     0;
     1878: diff =     0;
     1879: diff =     0;
     1880: diff =     0;
     1881: diff =     0;
     1882: diff =     0;
     1883: diff =     0;
     1884: diff =     0;
     1885: diff =     0;
     1886: diff =     0;
     1887: diff =     0;
     1888: diff =     0;
     1889: diff =     0;
     1890: diff =     0;
     1891: diff =     0;
     1892: diff =     0;
     1893: diff =     0;
     1894: diff =     0;
     1895: diff =     1;
     1896: diff =     1;
     1897: diff =     1;
     1898: diff =     1;
     1899: diff =     1;
     1900: diff =     1;
     1901: diff =     1;
     1902: diff =     1;
     1903: diff =     1;
     1904: diff =     1;
     1905: diff =     1;
     1906: diff =     1;
     1907: diff =     1;
     1908: diff =     1;
     1909: diff =     1;
     1910: diff =     1;
     1911: diff =     1;
     1912: diff =     1;
     1913: diff =     1;
     1914: diff =     1;
     1915: diff =     1;
     1916: diff =     1;
     1917: diff =     1;
     1918: diff =     1;
     1919: diff =     1;
     1920: diff =     0;
     1921: diff =     0;
     1922: diff =     0;
     1923: diff =     0;
     1924: diff =     0;
     1925: diff =     0;
     1926: diff =     0;
     1927: diff =     0;
     1928: diff =     0;
     1929: diff =     0;
     1930: diff =     0;
     1931: diff =     0;
     1932: diff =     0;
     1933: diff =     0;
     1934: diff =     0;
     1935: diff =     0;
     1936: diff =     0;
     1937: diff =     0;
     1938: diff =     0;
     1939: diff =     0;
     1940: diff =     0;
     1941: diff =     0;
     1942: diff =     0;
     1943: diff =     0;
     1944: diff =     0;
     1945: diff =     0;
     1946: diff =     0;
     1947: diff =     0;
     1948: diff =     0;
     1949: diff =     0;
     1950: diff =     0;
     1951: diff =     0;
     1952: diff =     0;
     1953: diff =     0;
     1954: diff =     0;
     1955: diff =     0;
     1956: diff =     0;
     1957: diff =     0;
     1958: diff =     0;
     1959: diff =     0;
     1960: diff =     0;
     1961: diff =     0;
     1962: diff =     0;
     1963: diff =     0;
     1964: diff =     0;
     1965: diff =     0;
     1966: diff =     0;
     1967: diff =     0;
     1968: diff =     0;
     1969: diff =     0;
     1970: diff =     0;
     1971: diff =     0;
     1972: diff =     0;
     1973: diff =     0;
     1974: diff =     0;
     1975: diff =     0;
     1976: diff =     0;
     1977: diff =     0;
     1978: diff =     0;
     1979: diff =     0;
     1980: diff =     0;
     1981: diff =     0;
     1982: diff =     0;
     1983: diff =     0;
     1984: diff =     0;
     1985: diff =     0;
     1986: diff =     0;
     1987: diff =     0;
     1988: diff =     0;
     1989: diff =     0;
     1990: diff =     0;
     1991: diff =     0;
     1992: diff =     0;
     1993: diff =     0;
     1994: diff =     0;
     1995: diff =     0;
     1996: diff =     0;
     1997: diff =     0;
     1998: diff =     0;
     1999: diff =     0;
     2000: diff =     0;
     2001: diff =     0;
     2002: diff =     0;
     2003: diff =     0;
     2004: diff =     0;
     2005: diff =     0;
     2006: diff =     0;
     2007: diff =     0;
     2008: diff =     0;
     2009: diff =     0;
     2010: diff =     0;
     2011: diff =     0;
     2012: diff =     0;
     2013: diff =     0;
     2014: diff =     0;
     2015: diff =     0;
     2016: diff =     0;
     2017: diff =     0;
     2018: diff =     0;
     2019: diff =     0;
     2020: diff =     0;
     2021: diff =     0;
     2022: diff =     0;
     2023: diff =     0;
     2024: diff =     0;
     2025: diff =     0;
     2026: diff =     1;
     2027: diff =     1;
     2028: diff =     1;
     2029: diff =     1;
     2030: diff =     1;
     2031: diff =     1;
     2032: diff =     1;
     2033: diff =     1;
     2034: diff =     1;
     2035: diff =     1;
     2036: diff =     1;
     2037: diff =     1;
     2038: diff =     1;
     2039: diff =     1;
     2040: diff =     1;
     2041: diff =     1;
     2042: diff =     1;
     2043: diff =     1;
     2044: diff =     1;
     2045: diff =     1;
     2046: diff =     1;
     2047: diff =     1;
    default: diff = 1;
    endcase
end
endmodule