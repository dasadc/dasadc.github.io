module sigmo_exact(output signed [13:0] y, input signed [11:0] x);
wire [11:0] xabs = (x>=0) ? x : -x;
reg signed [13:0] ytbl;
assign y = (x>=0) ? ytbl : 4096-ytbl;
always @* begin
    case (xabs)
    0: ytbl = 2048;
    1: ytbl = 2052;
    2: ytbl = 2056;
    3: ytbl = 2060;
    4: ytbl = 2064;
    5: ytbl = 2068;
    6: ytbl = 2072;
    7: ytbl = 2076;
    8: ytbl = 2080;
    9: ytbl = 2084;
    10: ytbl = 2088;
    11: ytbl = 2092;
    12: ytbl = 2096;
    13: ytbl = 2100;
    14: ytbl = 2104;
    15: ytbl = 2108;
    16: ytbl = 2112;
    17: ytbl = 2116;
    18: ytbl = 2120;
    19: ytbl = 2124;
    20: ytbl = 2128;
    21: ytbl = 2132;
    22: ytbl = 2136;
    23: ytbl = 2140;
    24: ytbl = 2144;
    25: ytbl = 2148;
    26: ytbl = 2152;
    27: ytbl = 2156;
    28: ytbl = 2160;
    29: ytbl = 2164;
    30: ytbl = 2168;
    31: ytbl = 2172;
    32: ytbl = 2176;
    33: ytbl = 2180;
    34: ytbl = 2184;
    35: ytbl = 2188;
    36: ytbl = 2192;
    37: ytbl = 2196;
    38: ytbl = 2200;
    39: ytbl = 2204;
    40: ytbl = 2208;
    41: ytbl = 2212;
    42: ytbl = 2216;
    43: ytbl = 2220;
    44: ytbl = 2224;
    45: ytbl = 2228;
    46: ytbl = 2232;
    47: ytbl = 2235;
    48: ytbl = 2239;
    49: ytbl = 2243;
    50: ytbl = 2247;
    51: ytbl = 2251;
    52: ytbl = 2255;
    53: ytbl = 2259;
    54: ytbl = 2263;
    55: ytbl = 2267;
    56: ytbl = 2271;
    57: ytbl = 2275;
    58: ytbl = 2279;
    59: ytbl = 2283;
    60: ytbl = 2287;
    61: ytbl = 2291;
    62: ytbl = 2295;
    63: ytbl = 2299;
    64: ytbl = 2303;
    65: ytbl = 2307;
    66: ytbl = 2311;
    67: ytbl = 2314;
    68: ytbl = 2318;
    69: ytbl = 2322;
    70: ytbl = 2326;
    71: ytbl = 2330;
    72: ytbl = 2334;
    73: ytbl = 2338;
    74: ytbl = 2342;
    75: ytbl = 2346;
    76: ytbl = 2350;
    77: ytbl = 2354;
    78: ytbl = 2358;
    79: ytbl = 2362;
    80: ytbl = 2365;
    81: ytbl = 2369;
    82: ytbl = 2373;
    83: ytbl = 2377;
    84: ytbl = 2381;
    85: ytbl = 2385;
    86: ytbl = 2389;
    87: ytbl = 2393;
    88: ytbl = 2397;
    89: ytbl = 2400;
    90: ytbl = 2404;
    91: ytbl = 2408;
    92: ytbl = 2412;
    93: ytbl = 2416;
    94: ytbl = 2420;
    95: ytbl = 2424;
    96: ytbl = 2428;
    97: ytbl = 2431;
    98: ytbl = 2435;
    99: ytbl = 2439;
    100: ytbl = 2443;
    101: ytbl = 2447;
    102: ytbl = 2451;
    103: ytbl = 2455;
    104: ytbl = 2458;
    105: ytbl = 2462;
    106: ytbl = 2466;
    107: ytbl = 2470;
    108: ytbl = 2474;
    109: ytbl = 2478;
    110: ytbl = 2481;
    111: ytbl = 2485;
    112: ytbl = 2489;
    113: ytbl = 2493;
    114: ytbl = 2497;
    115: ytbl = 2500;
    116: ytbl = 2504;
    117: ytbl = 2508;
    118: ytbl = 2512;
    119: ytbl = 2516;
    120: ytbl = 2519;
    121: ytbl = 2523;
    122: ytbl = 2527;
    123: ytbl = 2531;
    124: ytbl = 2535;
    125: ytbl = 2538;
    126: ytbl = 2542;
    127: ytbl = 2546;
    128: ytbl = 2550;
    129: ytbl = 2553;
    130: ytbl = 2557;
    131: ytbl = 2561;
    132: ytbl = 2565;
    133: ytbl = 2568;
    134: ytbl = 2572;
    135: ytbl = 2576;
    136: ytbl = 2580;
    137: ytbl = 2583;
    138: ytbl = 2587;
    139: ytbl = 2591;
    140: ytbl = 2594;
    141: ytbl = 2598;
    142: ytbl = 2602;
    143: ytbl = 2606;
    144: ytbl = 2609;
    145: ytbl = 2613;
    146: ytbl = 2617;
    147: ytbl = 2620;
    148: ytbl = 2624;
    149: ytbl = 2628;
    150: ytbl = 2631;
    151: ytbl = 2635;
    152: ytbl = 2639;
    153: ytbl = 2642;
    154: ytbl = 2646;
    155: ytbl = 2650;
    156: ytbl = 2653;
    157: ytbl = 2657;
    158: ytbl = 2661;
    159: ytbl = 2664;
    160: ytbl = 2668;
    161: ytbl = 2672;
    162: ytbl = 2675;
    163: ytbl = 2679;
    164: ytbl = 2682;
    165: ytbl = 2686;
    166: ytbl = 2690;
    167: ytbl = 2693;
    168: ytbl = 2697;
    169: ytbl = 2700;
    170: ytbl = 2704;
    171: ytbl = 2708;
    172: ytbl = 2711;
    173: ytbl = 2715;
    174: ytbl = 2718;
    175: ytbl = 2722;
    176: ytbl = 2726;
    177: ytbl = 2729;
    178: ytbl = 2733;
    179: ytbl = 2736;
    180: ytbl = 2740;
    181: ytbl = 2743;
    182: ytbl = 2747;
    183: ytbl = 2750;
    184: ytbl = 2754;
    185: ytbl = 2757;
    186: ytbl = 2761;
    187: ytbl = 2764;
    188: ytbl = 2768;
    189: ytbl = 2771;
    190: ytbl = 2775;
    191: ytbl = 2778;
    192: ytbl = 2782;
    193: ytbl = 2785;
    194: ytbl = 2789;
    195: ytbl = 2792;
    196: ytbl = 2796;
    197: ytbl = 2799;
    198: ytbl = 2803;
    199: ytbl = 2806;
    200: ytbl = 2810;
    201: ytbl = 2813;
    202: ytbl = 2817;
    203: ytbl = 2820;
    204: ytbl = 2823;
    205: ytbl = 2827;
    206: ytbl = 2830;
    207: ytbl = 2834;
    208: ytbl = 2837;
    209: ytbl = 2840;
    210: ytbl = 2844;
    211: ytbl = 2847;
    212: ytbl = 2851;
    213: ytbl = 2854;
    214: ytbl = 2857;
    215: ytbl = 2861;
    216: ytbl = 2864;
    217: ytbl = 2868;
    218: ytbl = 2871;
    219: ytbl = 2874;
    220: ytbl = 2878;
    221: ytbl = 2881;
    222: ytbl = 2884;
    223: ytbl = 2888;
    224: ytbl = 2891;
    225: ytbl = 2894;
    226: ytbl = 2898;
    227: ytbl = 2901;
    228: ytbl = 2904;
    229: ytbl = 2907;
    230: ytbl = 2911;
    231: ytbl = 2914;
    232: ytbl = 2917;
    233: ytbl = 2921;
    234: ytbl = 2924;
    235: ytbl = 2927;
    236: ytbl = 2930;
    237: ytbl = 2934;
    238: ytbl = 2937;
    239: ytbl = 2940;
    240: ytbl = 2943;
    241: ytbl = 2947;
    242: ytbl = 2950;
    243: ytbl = 2953;
    244: ytbl = 2956;
    245: ytbl = 2959;
    246: ytbl = 2963;
    247: ytbl = 2966;
    248: ytbl = 2969;
    249: ytbl = 2972;
    250: ytbl = 2975;
    251: ytbl = 2979;
    252: ytbl = 2982;
    253: ytbl = 2985;
    254: ytbl = 2988;
    255: ytbl = 2991;
    256: ytbl = 2994;
    257: ytbl = 2998;
    258: ytbl = 3001;
    259: ytbl = 3004;
    260: ytbl = 3007;
    261: ytbl = 3010;
    262: ytbl = 3013;
    263: ytbl = 3016;
    264: ytbl = 3019;
    265: ytbl = 3022;
    266: ytbl = 3026;
    267: ytbl = 3029;
    268: ytbl = 3032;
    269: ytbl = 3035;
    270: ytbl = 3038;
    271: ytbl = 3041;
    272: ytbl = 3044;
    273: ytbl = 3047;
    274: ytbl = 3050;
    275: ytbl = 3053;
    276: ytbl = 3056;
    277: ytbl = 3059;
    278: ytbl = 3062;
    279: ytbl = 3065;
    280: ytbl = 3068;
    281: ytbl = 3071;
    282: ytbl = 3074;
    283: ytbl = 3077;
    284: ytbl = 3080;
    285: ytbl = 3083;
    286: ytbl = 3086;
    287: ytbl = 3089;
    288: ytbl = 3092;
    289: ytbl = 3095;
    290: ytbl = 3098;
    291: ytbl = 3101;
    292: ytbl = 3104;
    293: ytbl = 3107;
    294: ytbl = 3110;
    295: ytbl = 3113;
    296: ytbl = 3116;
    297: ytbl = 3119;
    298: ytbl = 3121;
    299: ytbl = 3124;
    300: ytbl = 3127;
    301: ytbl = 3130;
    302: ytbl = 3133;
    303: ytbl = 3136;
    304: ytbl = 3139;
    305: ytbl = 3142;
    306: ytbl = 3144;
    307: ytbl = 3147;
    308: ytbl = 3150;
    309: ytbl = 3153;
    310: ytbl = 3156;
    311: ytbl = 3159;
    312: ytbl = 3161;
    313: ytbl = 3164;
    314: ytbl = 3167;
    315: ytbl = 3170;
    316: ytbl = 3173;
    317: ytbl = 3175;
    318: ytbl = 3178;
    319: ytbl = 3181;
    320: ytbl = 3184;
    321: ytbl = 3187;
    322: ytbl = 3189;
    323: ytbl = 3192;
    324: ytbl = 3195;
    325: ytbl = 3198;
    326: ytbl = 3200;
    327: ytbl = 3203;
    328: ytbl = 3206;
    329: ytbl = 3209;
    330: ytbl = 3211;
    331: ytbl = 3214;
    332: ytbl = 3217;
    333: ytbl = 3219;
    334: ytbl = 3222;
    335: ytbl = 3225;
    336: ytbl = 3227;
    337: ytbl = 3230;
    338: ytbl = 3233;
    339: ytbl = 3235;
    340: ytbl = 3238;
    341: ytbl = 3241;
    342: ytbl = 3243;
    343: ytbl = 3246;
    344: ytbl = 3249;
    345: ytbl = 3251;
    346: ytbl = 3254;
    347: ytbl = 3256;
    348: ytbl = 3259;
    349: ytbl = 3262;
    350: ytbl = 3264;
    351: ytbl = 3267;
    352: ytbl = 3269;
    353: ytbl = 3272;
    354: ytbl = 3275;
    355: ytbl = 3277;
    356: ytbl = 3280;
    357: ytbl = 3282;
    358: ytbl = 3285;
    359: ytbl = 3287;
    360: ytbl = 3290;
    361: ytbl = 3292;
    362: ytbl = 3295;
    363: ytbl = 3297;
    364: ytbl = 3300;
    365: ytbl = 3302;
    366: ytbl = 3305;
    367: ytbl = 3307;
    368: ytbl = 3310;
    369: ytbl = 3312;
    370: ytbl = 3315;
    371: ytbl = 3317;
    372: ytbl = 3320;
    373: ytbl = 3322;
    374: ytbl = 3325;
    375: ytbl = 3327;
    376: ytbl = 3330;
    377: ytbl = 3332;
    378: ytbl = 3334;
    379: ytbl = 3337;
    380: ytbl = 3339;
    381: ytbl = 3342;
    382: ytbl = 3344;
    383: ytbl = 3346;
    384: ytbl = 3349;
    385: ytbl = 3351;
    386: ytbl = 3354;
    387: ytbl = 3356;
    388: ytbl = 3358;
    389: ytbl = 3361;
    390: ytbl = 3363;
    391: ytbl = 3365;
    392: ytbl = 3368;
    393: ytbl = 3370;
    394: ytbl = 3372;
    395: ytbl = 3375;
    396: ytbl = 3377;
    397: ytbl = 3379;
    398: ytbl = 3382;
    399: ytbl = 3384;
    400: ytbl = 3386;
    401: ytbl = 3389;
    402: ytbl = 3391;
    403: ytbl = 3393;
    404: ytbl = 3395;
    405: ytbl = 3398;
    406: ytbl = 3400;
    407: ytbl = 3402;
    408: ytbl = 3404;
    409: ytbl = 3407;
    410: ytbl = 3409;
    411: ytbl = 3411;
    412: ytbl = 3413;
    413: ytbl = 3416;
    414: ytbl = 3418;
    415: ytbl = 3420;
    416: ytbl = 3422;
    417: ytbl = 3424;
    418: ytbl = 3427;
    419: ytbl = 3429;
    420: ytbl = 3431;
    421: ytbl = 3433;
    422: ytbl = 3435;
    423: ytbl = 3437;
    424: ytbl = 3440;
    425: ytbl = 3442;
    426: ytbl = 3444;
    427: ytbl = 3446;
    428: ytbl = 3448;
    429: ytbl = 3450;
    430: ytbl = 3452;
    431: ytbl = 3454;
    432: ytbl = 3457;
    433: ytbl = 3459;
    434: ytbl = 3461;
    435: ytbl = 3463;
    436: ytbl = 3465;
    437: ytbl = 3467;
    438: ytbl = 3469;
    439: ytbl = 3471;
    440: ytbl = 3473;
    441: ytbl = 3475;
    442: ytbl = 3477;
    443: ytbl = 3479;
    444: ytbl = 3481;
    445: ytbl = 3484;
    446: ytbl = 3486;
    447: ytbl = 3488;
    448: ytbl = 3490;
    449: ytbl = 3492;
    450: ytbl = 3494;
    451: ytbl = 3496;
    452: ytbl = 3498;
    453: ytbl = 3500;
    454: ytbl = 3502;
    455: ytbl = 3504;
    456: ytbl = 3506;
    457: ytbl = 3508;
    458: ytbl = 3510;
    459: ytbl = 3511;
    460: ytbl = 3513;
    461: ytbl = 3515;
    462: ytbl = 3517;
    463: ytbl = 3519;
    464: ytbl = 3521;
    465: ytbl = 3523;
    466: ytbl = 3525;
    467: ytbl = 3527;
    468: ytbl = 3529;
    469: ytbl = 3531;
    470: ytbl = 3533;
    471: ytbl = 3535;
    472: ytbl = 3536;
    473: ytbl = 3538;
    474: ytbl = 3540;
    475: ytbl = 3542;
    476: ytbl = 3544;
    477: ytbl = 3546;
    478: ytbl = 3548;
    479: ytbl = 3550;
    480: ytbl = 3551;
    481: ytbl = 3553;
    482: ytbl = 3555;
    483: ytbl = 3557;
    484: ytbl = 3559;
    485: ytbl = 3561;
    486: ytbl = 3562;
    487: ytbl = 3564;
    488: ytbl = 3566;
    489: ytbl = 3568;
    490: ytbl = 3570;
    491: ytbl = 3571;
    492: ytbl = 3573;
    493: ytbl = 3575;
    494: ytbl = 3577;
    495: ytbl = 3578;
    496: ytbl = 3580;
    497: ytbl = 3582;
    498: ytbl = 3584;
    499: ytbl = 3585;
    500: ytbl = 3587;
    501: ytbl = 3589;
    502: ytbl = 3591;
    503: ytbl = 3592;
    504: ytbl = 3594;
    505: ytbl = 3596;
    506: ytbl = 3598;
    507: ytbl = 3599;
    508: ytbl = 3601;
    509: ytbl = 3603;
    510: ytbl = 3604;
    511: ytbl = 3606;
    512: ytbl = 3608;
    513: ytbl = 3609;
    514: ytbl = 3611;
    515: ytbl = 3613;
    516: ytbl = 3614;
    517: ytbl = 3616;
    518: ytbl = 3618;
    519: ytbl = 3619;
    520: ytbl = 3621;
    521: ytbl = 3623;
    522: ytbl = 3624;
    523: ytbl = 3626;
    524: ytbl = 3628;
    525: ytbl = 3629;
    526: ytbl = 3631;
    527: ytbl = 3632;
    528: ytbl = 3634;
    529: ytbl = 3636;
    530: ytbl = 3637;
    531: ytbl = 3639;
    532: ytbl = 3640;
    533: ytbl = 3642;
    534: ytbl = 3644;
    535: ytbl = 3645;
    536: ytbl = 3647;
    537: ytbl = 3648;
    538: ytbl = 3650;
    539: ytbl = 3651;
    540: ytbl = 3653;
    541: ytbl = 3654;
    542: ytbl = 3656;
    543: ytbl = 3657;
    544: ytbl = 3659;
    545: ytbl = 3661;
    546: ytbl = 3662;
    547: ytbl = 3664;
    548: ytbl = 3665;
    549: ytbl = 3667;
    550: ytbl = 3668;
    551: ytbl = 3670;
    552: ytbl = 3671;
    553: ytbl = 3673;
    554: ytbl = 3674;
    555: ytbl = 3675;
    556: ytbl = 3677;
    557: ytbl = 3678;
    558: ytbl = 3680;
    559: ytbl = 3681;
    560: ytbl = 3683;
    561: ytbl = 3684;
    562: ytbl = 3686;
    563: ytbl = 3687;
    564: ytbl = 3689;
    565: ytbl = 3690;
    566: ytbl = 3691;
    567: ytbl = 3693;
    568: ytbl = 3694;
    569: ytbl = 3696;
    570: ytbl = 3697;
    571: ytbl = 3698;
    572: ytbl = 3700;
    573: ytbl = 3701;
    574: ytbl = 3703;
    575: ytbl = 3704;
    576: ytbl = 3705;
    577: ytbl = 3707;
    578: ytbl = 3708;
    579: ytbl = 3710;
    580: ytbl = 3711;
    581: ytbl = 3712;
    582: ytbl = 3714;
    583: ytbl = 3715;
    584: ytbl = 3716;
    585: ytbl = 3718;
    586: ytbl = 3719;
    587: ytbl = 3720;
    588: ytbl = 3722;
    589: ytbl = 3723;
    590: ytbl = 3724;
    591: ytbl = 3726;
    592: ytbl = 3727;
    593: ytbl = 3728;
    594: ytbl = 3730;
    595: ytbl = 3731;
    596: ytbl = 3732;
    597: ytbl = 3733;
    598: ytbl = 3735;
    599: ytbl = 3736;
    600: ytbl = 3737;
    601: ytbl = 3739;
    602: ytbl = 3740;
    603: ytbl = 3741;
    604: ytbl = 3742;
    605: ytbl = 3744;
    606: ytbl = 3745;
    607: ytbl = 3746;
    608: ytbl = 3747;
    609: ytbl = 3749;
    610: ytbl = 3750;
    611: ytbl = 3751;
    612: ytbl = 3752;
    613: ytbl = 3754;
    614: ytbl = 3755;
    615: ytbl = 3756;
    616: ytbl = 3757;
    617: ytbl = 3758;
    618: ytbl = 3760;
    619: ytbl = 3761;
    620: ytbl = 3762;
    621: ytbl = 3763;
    622: ytbl = 3764;
    623: ytbl = 3766;
    624: ytbl = 3767;
    625: ytbl = 3768;
    626: ytbl = 3769;
    627: ytbl = 3770;
    628: ytbl = 3772;
    629: ytbl = 3773;
    630: ytbl = 3774;
    631: ytbl = 3775;
    632: ytbl = 3776;
    633: ytbl = 3777;
    634: ytbl = 3778;
    635: ytbl = 3780;
    636: ytbl = 3781;
    637: ytbl = 3782;
    638: ytbl = 3783;
    639: ytbl = 3784;
    640: ytbl = 3785;
    641: ytbl = 3786;
    642: ytbl = 3788;
    643: ytbl = 3789;
    644: ytbl = 3790;
    645: ytbl = 3791;
    646: ytbl = 3792;
    647: ytbl = 3793;
    648: ytbl = 3794;
    649: ytbl = 3795;
    650: ytbl = 3796;
    651: ytbl = 3797;
    652: ytbl = 3798;
    653: ytbl = 3800;
    654: ytbl = 3801;
    655: ytbl = 3802;
    656: ytbl = 3803;
    657: ytbl = 3804;
    658: ytbl = 3805;
    659: ytbl = 3806;
    660: ytbl = 3807;
    661: ytbl = 3808;
    662: ytbl = 3809;
    663: ytbl = 3810;
    664: ytbl = 3811;
    665: ytbl = 3812;
    666: ytbl = 3813;
    667: ytbl = 3814;
    668: ytbl = 3815;
    669: ytbl = 3816;
    670: ytbl = 3817;
    671: ytbl = 3818;
    672: ytbl = 3819;
    673: ytbl = 3820;
    674: ytbl = 3821;
    675: ytbl = 3822;
    676: ytbl = 3823;
    677: ytbl = 3824;
    678: ytbl = 3825;
    679: ytbl = 3826;
    680: ytbl = 3827;
    681: ytbl = 3828;
    682: ytbl = 3829;
    683: ytbl = 3830;
    684: ytbl = 3831;
    685: ytbl = 3832;
    686: ytbl = 3833;
    687: ytbl = 3834;
    688: ytbl = 3835;
    689: ytbl = 3836;
    690: ytbl = 3837;
    691: ytbl = 3838;
    692: ytbl = 3839;
    693: ytbl = 3840;
    694: ytbl = 3841;
    695: ytbl = 3842;
    696: ytbl = 3843;
    697: ytbl = 3843;
    698: ytbl = 3844;
    699: ytbl = 3845;
    700: ytbl = 3846;
    701: ytbl = 3847;
    702: ytbl = 3848;
    703: ytbl = 3849;
    704: ytbl = 3850;
    705: ytbl = 3851;
    706: ytbl = 3852;
    707: ytbl = 3853;
    708: ytbl = 3853;
    709: ytbl = 3854;
    710: ytbl = 3855;
    711: ytbl = 3856;
    712: ytbl = 3857;
    713: ytbl = 3858;
    714: ytbl = 3859;
    715: ytbl = 3860;
    716: ytbl = 3861;
    717: ytbl = 3861;
    718: ytbl = 3862;
    719: ytbl = 3863;
    720: ytbl = 3864;
    721: ytbl = 3865;
    722: ytbl = 3866;
    723: ytbl = 3867;
    724: ytbl = 3867;
    725: ytbl = 3868;
    726: ytbl = 3869;
    727: ytbl = 3870;
    728: ytbl = 3871;
    729: ytbl = 3872;
    730: ytbl = 3872;
    731: ytbl = 3873;
    732: ytbl = 3874;
    733: ytbl = 3875;
    734: ytbl = 3876;
    735: ytbl = 3876;
    736: ytbl = 3877;
    737: ytbl = 3878;
    738: ytbl = 3879;
    739: ytbl = 3880;
    740: ytbl = 3880;
    741: ytbl = 3881;
    742: ytbl = 3882;
    743: ytbl = 3883;
    744: ytbl = 3884;
    745: ytbl = 3884;
    746: ytbl = 3885;
    747: ytbl = 3886;
    748: ytbl = 3887;
    749: ytbl = 3888;
    750: ytbl = 3888;
    751: ytbl = 3889;
    752: ytbl = 3890;
    753: ytbl = 3891;
    754: ytbl = 3891;
    755: ytbl = 3892;
    756: ytbl = 3893;
    757: ytbl = 3894;
    758: ytbl = 3894;
    759: ytbl = 3895;
    760: ytbl = 3896;
    761: ytbl = 3897;
    762: ytbl = 3897;
    763: ytbl = 3898;
    764: ytbl = 3899;
    765: ytbl = 3900;
    766: ytbl = 3900;
    767: ytbl = 3901;
    768: ytbl = 3902;
    769: ytbl = 3902;
    770: ytbl = 3903;
    771: ytbl = 3904;
    772: ytbl = 3905;
    773: ytbl = 3905;
    774: ytbl = 3906;
    775: ytbl = 3907;
    776: ytbl = 3907;
    777: ytbl = 3908;
    778: ytbl = 3909;
    779: ytbl = 3910;
    780: ytbl = 3910;
    781: ytbl = 3911;
    782: ytbl = 3912;
    783: ytbl = 3912;
    784: ytbl = 3913;
    785: ytbl = 3914;
    786: ytbl = 3914;
    787: ytbl = 3915;
    788: ytbl = 3916;
    789: ytbl = 3916;
    790: ytbl = 3917;
    791: ytbl = 3918;
    792: ytbl = 3918;
    793: ytbl = 3919;
    794: ytbl = 3920;
    795: ytbl = 3920;
    796: ytbl = 3921;
    797: ytbl = 3922;
    798: ytbl = 3922;
    799: ytbl = 3923;
    800: ytbl = 3924;
    801: ytbl = 3924;
    802: ytbl = 3925;
    803: ytbl = 3926;
    804: ytbl = 3926;
    805: ytbl = 3927;
    806: ytbl = 3927;
    807: ytbl = 3928;
    808: ytbl = 3929;
    809: ytbl = 3929;
    810: ytbl = 3930;
    811: ytbl = 3931;
    812: ytbl = 3931;
    813: ytbl = 3932;
    814: ytbl = 3932;
    815: ytbl = 3933;
    816: ytbl = 3934;
    817: ytbl = 3934;
    818: ytbl = 3935;
    819: ytbl = 3935;
    820: ytbl = 3936;
    821: ytbl = 3937;
    822: ytbl = 3937;
    823: ytbl = 3938;
    824: ytbl = 3938;
    825: ytbl = 3939;
    826: ytbl = 3940;
    827: ytbl = 3940;
    828: ytbl = 3941;
    829: ytbl = 3941;
    830: ytbl = 3942;
    831: ytbl = 3943;
    832: ytbl = 3943;
    833: ytbl = 3944;
    834: ytbl = 3944;
    835: ytbl = 3945;
    836: ytbl = 3945;
    837: ytbl = 3946;
    838: ytbl = 3947;
    839: ytbl = 3947;
    840: ytbl = 3948;
    841: ytbl = 3948;
    842: ytbl = 3949;
    843: ytbl = 3949;
    844: ytbl = 3950;
    845: ytbl = 3950;
    846: ytbl = 3951;
    847: ytbl = 3952;
    848: ytbl = 3952;
    849: ytbl = 3953;
    850: ytbl = 3953;
    851: ytbl = 3954;
    852: ytbl = 3954;
    853: ytbl = 3955;
    854: ytbl = 3955;
    855: ytbl = 3956;
    856: ytbl = 3956;
    857: ytbl = 3957;
    858: ytbl = 3957;
    859: ytbl = 3958;
    860: ytbl = 3958;
    861: ytbl = 3959;
    862: ytbl = 3959;
    863: ytbl = 3960;
    864: ytbl = 3960;
    865: ytbl = 3961;
    866: ytbl = 3961;
    867: ytbl = 3962;
    868: ytbl = 3963;
    869: ytbl = 3963;
    870: ytbl = 3964;
    871: ytbl = 3964;
    872: ytbl = 3965;
    873: ytbl = 3965;
    874: ytbl = 3966;
    875: ytbl = 3966;
    876: ytbl = 3966;
    877: ytbl = 3967;
    878: ytbl = 3967;
    879: ytbl = 3968;
    880: ytbl = 3968;
    881: ytbl = 3969;
    882: ytbl = 3969;
    883: ytbl = 3970;
    884: ytbl = 3970;
    885: ytbl = 3971;
    886: ytbl = 3971;
    887: ytbl = 3972;
    888: ytbl = 3972;
    889: ytbl = 3973;
    890: ytbl = 3973;
    891: ytbl = 3974;
    892: ytbl = 3974;
    893: ytbl = 3975;
    894: ytbl = 3975;
    895: ytbl = 3975;
    896: ytbl = 3976;
    897: ytbl = 3976;
    898: ytbl = 3977;
    899: ytbl = 3977;
    900: ytbl = 3978;
    901: ytbl = 3978;
    902: ytbl = 3979;
    903: ytbl = 3979;
    904: ytbl = 3980;
    905: ytbl = 3980;
    906: ytbl = 3980;
    907: ytbl = 3981;
    908: ytbl = 3981;
    909: ytbl = 3982;
    910: ytbl = 3982;
    911: ytbl = 3983;
    912: ytbl = 3983;
    913: ytbl = 3983;
    914: ytbl = 3984;
    915: ytbl = 3984;
    916: ytbl = 3985;
    917: ytbl = 3985;
    918: ytbl = 3986;
    919: ytbl = 3986;
    920: ytbl = 3986;
    921: ytbl = 3987;
    922: ytbl = 3987;
    923: ytbl = 3988;
    924: ytbl = 3988;
    925: ytbl = 3988;
    926: ytbl = 3989;
    927: ytbl = 3989;
    928: ytbl = 3990;
    929: ytbl = 3990;
    930: ytbl = 3990;
    931: ytbl = 3991;
    932: ytbl = 3991;
    933: ytbl = 3992;
    934: ytbl = 3992;
    935: ytbl = 3992;
    936: ytbl = 3993;
    937: ytbl = 3993;
    938: ytbl = 3994;
    939: ytbl = 3994;
    940: ytbl = 3994;
    941: ytbl = 3995;
    942: ytbl = 3995;
    943: ytbl = 3996;
    944: ytbl = 3996;
    945: ytbl = 3996;
    946: ytbl = 3997;
    947: ytbl = 3997;
    948: ytbl = 3997;
    949: ytbl = 3998;
    950: ytbl = 3998;
    951: ytbl = 3999;
    952: ytbl = 3999;
    953: ytbl = 3999;
    954: ytbl = 4000;
    955: ytbl = 4000;
    956: ytbl = 4000;
    957: ytbl = 4001;
    958: ytbl = 4001;
    959: ytbl = 4002;
    960: ytbl = 4002;
    961: ytbl = 4002;
    962: ytbl = 4003;
    963: ytbl = 4003;
    964: ytbl = 4003;
    965: ytbl = 4004;
    966: ytbl = 4004;
    967: ytbl = 4004;
    968: ytbl = 4005;
    969: ytbl = 4005;
    970: ytbl = 4005;
    971: ytbl = 4006;
    972: ytbl = 4006;
    973: ytbl = 4006;
    974: ytbl = 4007;
    975: ytbl = 4007;
    976: ytbl = 4007;
    977: ytbl = 4008;
    978: ytbl = 4008;
    979: ytbl = 4008;
    980: ytbl = 4009;
    981: ytbl = 4009;
    982: ytbl = 4009;
    983: ytbl = 4010;
    984: ytbl = 4010;
    985: ytbl = 4010;
    986: ytbl = 4011;
    987: ytbl = 4011;
    988: ytbl = 4011;
    989: ytbl = 4012;
    990: ytbl = 4012;
    991: ytbl = 4012;
    992: ytbl = 4013;
    993: ytbl = 4013;
    994: ytbl = 4013;
    995: ytbl = 4014;
    996: ytbl = 4014;
    997: ytbl = 4014;
    998: ytbl = 4015;
    999: ytbl = 4015;
    1000: ytbl = 4015;
    1001: ytbl = 4016;
    1002: ytbl = 4016;
    1003: ytbl = 4016;
    1004: ytbl = 4016;
    1005: ytbl = 4017;
    1006: ytbl = 4017;
    1007: ytbl = 4017;
    1008: ytbl = 4018;
    1009: ytbl = 4018;
    1010: ytbl = 4018;
    1011: ytbl = 4019;
    1012: ytbl = 4019;
    1013: ytbl = 4019;
    1014: ytbl = 4019;
    1015: ytbl = 4020;
    1016: ytbl = 4020;
    1017: ytbl = 4020;
    1018: ytbl = 4021;
    1019: ytbl = 4021;
    1020: ytbl = 4021;
    1021: ytbl = 4021;
    1022: ytbl = 4022;
    1023: ytbl = 4022;
    1024: ytbl = 4022;
    1025: ytbl = 4023;
    1026: ytbl = 4023;
    1027: ytbl = 4023;
    1028: ytbl = 4023;
    1029: ytbl = 4024;
    1030: ytbl = 4024;
    1031: ytbl = 4024;
    1032: ytbl = 4025;
    1033: ytbl = 4025;
    1034: ytbl = 4025;
    1035: ytbl = 4025;
    1036: ytbl = 4026;
    1037: ytbl = 4026;
    1038: ytbl = 4026;
    1039: ytbl = 4026;
    1040: ytbl = 4027;
    1041: ytbl = 4027;
    1042: ytbl = 4027;
    1043: ytbl = 4028;
    1044: ytbl = 4028;
    1045: ytbl = 4028;
    1046: ytbl = 4028;
    1047: ytbl = 4029;
    1048: ytbl = 4029;
    1049: ytbl = 4029;
    1050: ytbl = 4029;
    1051: ytbl = 4030;
    1052: ytbl = 4030;
    1053: ytbl = 4030;
    1054: ytbl = 4030;
    1055: ytbl = 4031;
    1056: ytbl = 4031;
    1057: ytbl = 4031;
    1058: ytbl = 4031;
    1059: ytbl = 4032;
    1060: ytbl = 4032;
    1061: ytbl = 4032;
    1062: ytbl = 4032;
    1063: ytbl = 4033;
    1064: ytbl = 4033;
    1065: ytbl = 4033;
    1066: ytbl = 4033;
    1067: ytbl = 4034;
    1068: ytbl = 4034;
    1069: ytbl = 4034;
    1070: ytbl = 4034;
    1071: ytbl = 4034;
    1072: ytbl = 4035;
    1073: ytbl = 4035;
    1074: ytbl = 4035;
    1075: ytbl = 4035;
    1076: ytbl = 4036;
    1077: ytbl = 4036;
    1078: ytbl = 4036;
    1079: ytbl = 4036;
    1080: ytbl = 4037;
    1081: ytbl = 4037;
    1082: ytbl = 4037;
    1083: ytbl = 4037;
    1084: ytbl = 4038;
    1085: ytbl = 4038;
    1086: ytbl = 4038;
    1087: ytbl = 4038;
    1088: ytbl = 4038;
    1089: ytbl = 4039;
    1090: ytbl = 4039;
    1091: ytbl = 4039;
    1092: ytbl = 4039;
    1093: ytbl = 4039;
    1094: ytbl = 4040;
    1095: ytbl = 4040;
    1096: ytbl = 4040;
    1097: ytbl = 4040;
    1098: ytbl = 4041;
    1099: ytbl = 4041;
    1100: ytbl = 4041;
    1101: ytbl = 4041;
    1102: ytbl = 4041;
    1103: ytbl = 4042;
    1104: ytbl = 4042;
    1105: ytbl = 4042;
    1106: ytbl = 4042;
    1107: ytbl = 4042;
    1108: ytbl = 4043;
    1109: ytbl = 4043;
    1110: ytbl = 4043;
    1111: ytbl = 4043;
    1112: ytbl = 4043;
    1113: ytbl = 4044;
    1114: ytbl = 4044;
    1115: ytbl = 4044;
    1116: ytbl = 4044;
    1117: ytbl = 4044;
    1118: ytbl = 4045;
    1119: ytbl = 4045;
    1120: ytbl = 4045;
    1121: ytbl = 4045;
    1122: ytbl = 4045;
    1123: ytbl = 4046;
    1124: ytbl = 4046;
    1125: ytbl = 4046;
    1126: ytbl = 4046;
    1127: ytbl = 4046;
    1128: ytbl = 4047;
    1129: ytbl = 4047;
    1130: ytbl = 4047;
    1131: ytbl = 4047;
    1132: ytbl = 4047;
    1133: ytbl = 4048;
    1134: ytbl = 4048;
    1135: ytbl = 4048;
    1136: ytbl = 4048;
    1137: ytbl = 4048;
    1138: ytbl = 4048;
    1139: ytbl = 4049;
    1140: ytbl = 4049;
    1141: ytbl = 4049;
    1142: ytbl = 4049;
    1143: ytbl = 4049;
    1144: ytbl = 4050;
    1145: ytbl = 4050;
    1146: ytbl = 4050;
    1147: ytbl = 4050;
    1148: ytbl = 4050;
    1149: ytbl = 4050;
    1150: ytbl = 4051;
    1151: ytbl = 4051;
    1152: ytbl = 4051;
    1153: ytbl = 4051;
    1154: ytbl = 4051;
    1155: ytbl = 4052;
    1156: ytbl = 4052;
    1157: ytbl = 4052;
    1158: ytbl = 4052;
    1159: ytbl = 4052;
    1160: ytbl = 4052;
    1161: ytbl = 4053;
    1162: ytbl = 4053;
    1163: ytbl = 4053;
    1164: ytbl = 4053;
    1165: ytbl = 4053;
    1166: ytbl = 4053;
    1167: ytbl = 4054;
    1168: ytbl = 4054;
    1169: ytbl = 4054;
    1170: ytbl = 4054;
    1171: ytbl = 4054;
    1172: ytbl = 4054;
    1173: ytbl = 4055;
    1174: ytbl = 4055;
    1175: ytbl = 4055;
    1176: ytbl = 4055;
    1177: ytbl = 4055;
    1178: ytbl = 4055;
    1179: ytbl = 4055;
    1180: ytbl = 4056;
    1181: ytbl = 4056;
    1182: ytbl = 4056;
    1183: ytbl = 4056;
    1184: ytbl = 4056;
    1185: ytbl = 4056;
    1186: ytbl = 4057;
    1187: ytbl = 4057;
    1188: ytbl = 4057;
    1189: ytbl = 4057;
    1190: ytbl = 4057;
    1191: ytbl = 4057;
    1192: ytbl = 4057;
    1193: ytbl = 4058;
    1194: ytbl = 4058;
    1195: ytbl = 4058;
    1196: ytbl = 4058;
    1197: ytbl = 4058;
    1198: ytbl = 4058;
    1199: ytbl = 4058;
    1200: ytbl = 4059;
    1201: ytbl = 4059;
    1202: ytbl = 4059;
    1203: ytbl = 4059;
    1204: ytbl = 4059;
    1205: ytbl = 4059;
    1206: ytbl = 4059;
    1207: ytbl = 4060;
    1208: ytbl = 4060;
    1209: ytbl = 4060;
    1210: ytbl = 4060;
    1211: ytbl = 4060;
    1212: ytbl = 4060;
    1213: ytbl = 4060;
    1214: ytbl = 4061;
    1215: ytbl = 4061;
    1216: ytbl = 4061;
    1217: ytbl = 4061;
    1218: ytbl = 4061;
    1219: ytbl = 4061;
    1220: ytbl = 4061;
    1221: ytbl = 4062;
    1222: ytbl = 4062;
    1223: ytbl = 4062;
    1224: ytbl = 4062;
    1225: ytbl = 4062;
    1226: ytbl = 4062;
    1227: ytbl = 4062;
    1228: ytbl = 4062;
    1229: ytbl = 4063;
    1230: ytbl = 4063;
    1231: ytbl = 4063;
    1232: ytbl = 4063;
    1233: ytbl = 4063;
    1234: ytbl = 4063;
    1235: ytbl = 4063;
    1236: ytbl = 4063;
    1237: ytbl = 4064;
    1238: ytbl = 4064;
    1239: ytbl = 4064;
    1240: ytbl = 4064;
    1241: ytbl = 4064;
    1242: ytbl = 4064;
    1243: ytbl = 4064;
    1244: ytbl = 4064;
    1245: ytbl = 4065;
    1246: ytbl = 4065;
    1247: ytbl = 4065;
    1248: ytbl = 4065;
    1249: ytbl = 4065;
    1250: ytbl = 4065;
    1251: ytbl = 4065;
    1252: ytbl = 4065;
    1253: ytbl = 4066;
    1254: ytbl = 4066;
    1255: ytbl = 4066;
    1256: ytbl = 4066;
    1257: ytbl = 4066;
    1258: ytbl = 4066;
    1259: ytbl = 4066;
    1260: ytbl = 4066;
    1261: ytbl = 4066;
    1262: ytbl = 4067;
    1263: ytbl = 4067;
    1264: ytbl = 4067;
    1265: ytbl = 4067;
    1266: ytbl = 4067;
    1267: ytbl = 4067;
    1268: ytbl = 4067;
    1269: ytbl = 4067;
    1270: ytbl = 4068;
    1271: ytbl = 4068;
    1272: ytbl = 4068;
    1273: ytbl = 4068;
    1274: ytbl = 4068;
    1275: ytbl = 4068;
    1276: ytbl = 4068;
    1277: ytbl = 4068;
    1278: ytbl = 4068;
    1279: ytbl = 4068;
    1280: ytbl = 4069;
    1281: ytbl = 4069;
    1282: ytbl = 4069;
    1283: ytbl = 4069;
    1284: ytbl = 4069;
    1285: ytbl = 4069;
    1286: ytbl = 4069;
    1287: ytbl = 4069;
    1288: ytbl = 4069;
    1289: ytbl = 4070;
    1290: ytbl = 4070;
    1291: ytbl = 4070;
    1292: ytbl = 4070;
    1293: ytbl = 4070;
    1294: ytbl = 4070;
    1295: ytbl = 4070;
    1296: ytbl = 4070;
    1297: ytbl = 4070;
    1298: ytbl = 4070;
    1299: ytbl = 4071;
    1300: ytbl = 4071;
    1301: ytbl = 4071;
    1302: ytbl = 4071;
    1303: ytbl = 4071;
    1304: ytbl = 4071;
    1305: ytbl = 4071;
    1306: ytbl = 4071;
    1307: ytbl = 4071;
    1308: ytbl = 4071;
    1309: ytbl = 4072;
    1310: ytbl = 4072;
    1311: ytbl = 4072;
    1312: ytbl = 4072;
    1313: ytbl = 4072;
    1314: ytbl = 4072;
    1315: ytbl = 4072;
    1316: ytbl = 4072;
    1317: ytbl = 4072;
    1318: ytbl = 4072;
    1319: ytbl = 4072;
    1320: ytbl = 4073;
    1321: ytbl = 4073;
    1322: ytbl = 4073;
    1323: ytbl = 4073;
    1324: ytbl = 4073;
    1325: ytbl = 4073;
    1326: ytbl = 4073;
    1327: ytbl = 4073;
    1328: ytbl = 4073;
    1329: ytbl = 4073;
    1330: ytbl = 4073;
    1331: ytbl = 4074;
    1332: ytbl = 4074;
    1333: ytbl = 4074;
    1334: ytbl = 4074;
    1335: ytbl = 4074;
    1336: ytbl = 4074;
    1337: ytbl = 4074;
    1338: ytbl = 4074;
    1339: ytbl = 4074;
    1340: ytbl = 4074;
    1341: ytbl = 4074;
    1342: ytbl = 4074;
    1343: ytbl = 4075;
    1344: ytbl = 4075;
    1345: ytbl = 4075;
    1346: ytbl = 4075;
    1347: ytbl = 4075;
    1348: ytbl = 4075;
    1349: ytbl = 4075;
    1350: ytbl = 4075;
    1351: ytbl = 4075;
    1352: ytbl = 4075;
    1353: ytbl = 4075;
    1354: ytbl = 4075;
    1355: ytbl = 4076;
    1356: ytbl = 4076;
    1357: ytbl = 4076;
    1358: ytbl = 4076;
    1359: ytbl = 4076;
    1360: ytbl = 4076;
    1361: ytbl = 4076;
    1362: ytbl = 4076;
    1363: ytbl = 4076;
    1364: ytbl = 4076;
    1365: ytbl = 4076;
    1366: ytbl = 4076;
    1367: ytbl = 4076;
    1368: ytbl = 4077;
    1369: ytbl = 4077;
    1370: ytbl = 4077;
    1371: ytbl = 4077;
    1372: ytbl = 4077;
    1373: ytbl = 4077;
    1374: ytbl = 4077;
    1375: ytbl = 4077;
    1376: ytbl = 4077;
    1377: ytbl = 4077;
    1378: ytbl = 4077;
    1379: ytbl = 4077;
    1380: ytbl = 4077;
    1381: ytbl = 4077;
    1382: ytbl = 4078;
    1383: ytbl = 4078;
    1384: ytbl = 4078;
    1385: ytbl = 4078;
    1386: ytbl = 4078;
    1387: ytbl = 4078;
    1388: ytbl = 4078;
    1389: ytbl = 4078;
    1390: ytbl = 4078;
    1391: ytbl = 4078;
    1392: ytbl = 4078;
    1393: ytbl = 4078;
    1394: ytbl = 4078;
    1395: ytbl = 4078;
    1396: ytbl = 4079;
    1397: ytbl = 4079;
    1398: ytbl = 4079;
    1399: ytbl = 4079;
    1400: ytbl = 4079;
    1401: ytbl = 4079;
    1402: ytbl = 4079;
    1403: ytbl = 4079;
    1404: ytbl = 4079;
    1405: ytbl = 4079;
    1406: ytbl = 4079;
    1407: ytbl = 4079;
    1408: ytbl = 4079;
    1409: ytbl = 4079;
    1410: ytbl = 4079;
    1411: ytbl = 4080;
    1412: ytbl = 4080;
    1413: ytbl = 4080;
    1414: ytbl = 4080;
    1415: ytbl = 4080;
    1416: ytbl = 4080;
    1417: ytbl = 4080;
    1418: ytbl = 4080;
    1419: ytbl = 4080;
    1420: ytbl = 4080;
    1421: ytbl = 4080;
    1422: ytbl = 4080;
    1423: ytbl = 4080;
    1424: ytbl = 4080;
    1425: ytbl = 4080;
    1426: ytbl = 4080;
    1427: ytbl = 4081;
    1428: ytbl = 4081;
    1429: ytbl = 4081;
    1430: ytbl = 4081;
    1431: ytbl = 4081;
    1432: ytbl = 4081;
    1433: ytbl = 4081;
    1434: ytbl = 4081;
    1435: ytbl = 4081;
    1436: ytbl = 4081;
    1437: ytbl = 4081;
    1438: ytbl = 4081;
    1439: ytbl = 4081;
    1440: ytbl = 4081;
    1441: ytbl = 4081;
    1442: ytbl = 4081;
    1443: ytbl = 4081;
    1444: ytbl = 4082;
    1445: ytbl = 4082;
    1446: ytbl = 4082;
    1447: ytbl = 4082;
    1448: ytbl = 4082;
    1449: ytbl = 4082;
    1450: ytbl = 4082;
    1451: ytbl = 4082;
    1452: ytbl = 4082;
    1453: ytbl = 4082;
    1454: ytbl = 4082;
    1455: ytbl = 4082;
    1456: ytbl = 4082;
    1457: ytbl = 4082;
    1458: ytbl = 4082;
    1459: ytbl = 4082;
    1460: ytbl = 4082;
    1461: ytbl = 4082;
    1462: ytbl = 4082;
    1463: ytbl = 4083;
    1464: ytbl = 4083;
    1465: ytbl = 4083;
    1466: ytbl = 4083;
    1467: ytbl = 4083;
    1468: ytbl = 4083;
    1469: ytbl = 4083;
    1470: ytbl = 4083;
    1471: ytbl = 4083;
    1472: ytbl = 4083;
    1473: ytbl = 4083;
    1474: ytbl = 4083;
    1475: ytbl = 4083;
    1476: ytbl = 4083;
    1477: ytbl = 4083;
    1478: ytbl = 4083;
    1479: ytbl = 4083;
    1480: ytbl = 4083;
    1481: ytbl = 4083;
    1482: ytbl = 4084;
    1483: ytbl = 4084;
    1484: ytbl = 4084;
    1485: ytbl = 4084;
    1486: ytbl = 4084;
    1487: ytbl = 4084;
    1488: ytbl = 4084;
    1489: ytbl = 4084;
    1490: ytbl = 4084;
    1491: ytbl = 4084;
    1492: ytbl = 4084;
    1493: ytbl = 4084;
    1494: ytbl = 4084;
    1495: ytbl = 4084;
    1496: ytbl = 4084;
    1497: ytbl = 4084;
    1498: ytbl = 4084;
    1499: ytbl = 4084;
    1500: ytbl = 4084;
    1501: ytbl = 4084;
    1502: ytbl = 4084;
    1503: ytbl = 4084;
    1504: ytbl = 4085;
    1505: ytbl = 4085;
    1506: ytbl = 4085;
    1507: ytbl = 4085;
    1508: ytbl = 4085;
    1509: ytbl = 4085;
    1510: ytbl = 4085;
    1511: ytbl = 4085;
    1512: ytbl = 4085;
    1513: ytbl = 4085;
    1514: ytbl = 4085;
    1515: ytbl = 4085;
    1516: ytbl = 4085;
    1517: ytbl = 4085;
    1518: ytbl = 4085;
    1519: ytbl = 4085;
    1520: ytbl = 4085;
    1521: ytbl = 4085;
    1522: ytbl = 4085;
    1523: ytbl = 4085;
    1524: ytbl = 4085;
    1525: ytbl = 4085;
    1526: ytbl = 4085;
    1527: ytbl = 4086;
    1528: ytbl = 4086;
    1529: ytbl = 4086;
    1530: ytbl = 4086;
    1531: ytbl = 4086;
    1532: ytbl = 4086;
    1533: ytbl = 4086;
    1534: ytbl = 4086;
    1535: ytbl = 4086;
    1536: ytbl = 4086;
    1537: ytbl = 4086;
    1538: ytbl = 4086;
    1539: ytbl = 4086;
    1540: ytbl = 4086;
    1541: ytbl = 4086;
    1542: ytbl = 4086;
    1543: ytbl = 4086;
    1544: ytbl = 4086;
    1545: ytbl = 4086;
    1546: ytbl = 4086;
    1547: ytbl = 4086;
    1548: ytbl = 4086;
    1549: ytbl = 4086;
    1550: ytbl = 4086;
    1551: ytbl = 4086;
    1552: ytbl = 4086;
    1553: ytbl = 4087;
    1554: ytbl = 4087;
    1555: ytbl = 4087;
    1556: ytbl = 4087;
    1557: ytbl = 4087;
    1558: ytbl = 4087;
    1559: ytbl = 4087;
    1560: ytbl = 4087;
    1561: ytbl = 4087;
    1562: ytbl = 4087;
    1563: ytbl = 4087;
    1564: ytbl = 4087;
    1565: ytbl = 4087;
    1566: ytbl = 4087;
    1567: ytbl = 4087;
    1568: ytbl = 4087;
    1569: ytbl = 4087;
    1570: ytbl = 4087;
    1571: ytbl = 4087;
    1572: ytbl = 4087;
    1573: ytbl = 4087;
    1574: ytbl = 4087;
    1575: ytbl = 4087;
    1576: ytbl = 4087;
    1577: ytbl = 4087;
    1578: ytbl = 4087;
    1579: ytbl = 4087;
    1580: ytbl = 4087;
    1581: ytbl = 4088;
    1582: ytbl = 4088;
    1583: ytbl = 4088;
    1584: ytbl = 4088;
    1585: ytbl = 4088;
    1586: ytbl = 4088;
    1587: ytbl = 4088;
    1588: ytbl = 4088;
    1589: ytbl = 4088;
    1590: ytbl = 4088;
    1591: ytbl = 4088;
    1592: ytbl = 4088;
    1593: ytbl = 4088;
    1594: ytbl = 4088;
    1595: ytbl = 4088;
    1596: ytbl = 4088;
    1597: ytbl = 4088;
    1598: ytbl = 4088;
    1599: ytbl = 4088;
    1600: ytbl = 4088;
    1601: ytbl = 4088;
    1602: ytbl = 4088;
    1603: ytbl = 4088;
    1604: ytbl = 4088;
    1605: ytbl = 4088;
    1606: ytbl = 4088;
    1607: ytbl = 4088;
    1608: ytbl = 4088;
    1609: ytbl = 4088;
    1610: ytbl = 4088;
    1611: ytbl = 4088;
    1612: ytbl = 4088;
    1613: ytbl = 4088;
    1614: ytbl = 4089;
    1615: ytbl = 4089;
    1616: ytbl = 4089;
    1617: ytbl = 4089;
    1618: ytbl = 4089;
    1619: ytbl = 4089;
    1620: ytbl = 4089;
    1621: ytbl = 4089;
    1622: ytbl = 4089;
    1623: ytbl = 4089;
    1624: ytbl = 4089;
    1625: ytbl = 4089;
    1626: ytbl = 4089;
    1627: ytbl = 4089;
    1628: ytbl = 4089;
    1629: ytbl = 4089;
    1630: ytbl = 4089;
    1631: ytbl = 4089;
    1632: ytbl = 4089;
    1633: ytbl = 4089;
    1634: ytbl = 4089;
    1635: ytbl = 4089;
    1636: ytbl = 4089;
    1637: ytbl = 4089;
    1638: ytbl = 4089;
    1639: ytbl = 4089;
    1640: ytbl = 4089;
    1641: ytbl = 4089;
    1642: ytbl = 4089;
    1643: ytbl = 4089;
    1644: ytbl = 4089;
    1645: ytbl = 4089;
    1646: ytbl = 4089;
    1647: ytbl = 4089;
    1648: ytbl = 4089;
    1649: ytbl = 4089;
    1650: ytbl = 4090;
    1651: ytbl = 4090;
    1652: ytbl = 4090;
    1653: ytbl = 4090;
    1654: ytbl = 4090;
    1655: ytbl = 4090;
    1656: ytbl = 4090;
    1657: ytbl = 4090;
    1658: ytbl = 4090;
    1659: ytbl = 4090;
    1660: ytbl = 4090;
    1661: ytbl = 4090;
    1662: ytbl = 4090;
    1663: ytbl = 4090;
    1664: ytbl = 4090;
    1665: ytbl = 4090;
    1666: ytbl = 4090;
    1667: ytbl = 4090;
    1668: ytbl = 4090;
    1669: ytbl = 4090;
    1670: ytbl = 4090;
    1671: ytbl = 4090;
    1672: ytbl = 4090;
    1673: ytbl = 4090;
    1674: ytbl = 4090;
    1675: ytbl = 4090;
    1676: ytbl = 4090;
    1677: ytbl = 4090;
    1678: ytbl = 4090;
    1679: ytbl = 4090;
    1680: ytbl = 4090;
    1681: ytbl = 4090;
    1682: ytbl = 4090;
    1683: ytbl = 4090;
    1684: ytbl = 4090;
    1685: ytbl = 4090;
    1686: ytbl = 4090;
    1687: ytbl = 4090;
    1688: ytbl = 4090;
    1689: ytbl = 4090;
    1690: ytbl = 4090;
    1691: ytbl = 4090;
    1692: ytbl = 4090;
    1693: ytbl = 4091;
    1694: ytbl = 4091;
    1695: ytbl = 4091;
    1696: ytbl = 4091;
    1697: ytbl = 4091;
    1698: ytbl = 4091;
    1699: ytbl = 4091;
    1700: ytbl = 4091;
    1701: ytbl = 4091;
    1702: ytbl = 4091;
    1703: ytbl = 4091;
    1704: ytbl = 4091;
    1705: ytbl = 4091;
    1706: ytbl = 4091;
    1707: ytbl = 4091;
    1708: ytbl = 4091;
    1709: ytbl = 4091;
    1710: ytbl = 4091;
    1711: ytbl = 4091;
    1712: ytbl = 4091;
    1713: ytbl = 4091;
    1714: ytbl = 4091;
    1715: ytbl = 4091;
    1716: ytbl = 4091;
    1717: ytbl = 4091;
    1718: ytbl = 4091;
    1719: ytbl = 4091;
    1720: ytbl = 4091;
    1721: ytbl = 4091;
    1722: ytbl = 4091;
    1723: ytbl = 4091;
    1724: ytbl = 4091;
    1725: ytbl = 4091;
    1726: ytbl = 4091;
    1727: ytbl = 4091;
    1728: ytbl = 4091;
    1729: ytbl = 4091;
    1730: ytbl = 4091;
    1731: ytbl = 4091;
    1732: ytbl = 4091;
    1733: ytbl = 4091;
    1734: ytbl = 4091;
    1735: ytbl = 4091;
    1736: ytbl = 4091;
    1737: ytbl = 4091;
    1738: ytbl = 4091;
    1739: ytbl = 4091;
    1740: ytbl = 4091;
    1741: ytbl = 4091;
    1742: ytbl = 4091;
    1743: ytbl = 4091;
    1744: ytbl = 4091;
    1745: ytbl = 4092;
    1746: ytbl = 4092;
    1747: ytbl = 4092;
    1748: ytbl = 4092;
    1749: ytbl = 4092;
    1750: ytbl = 4092;
    1751: ytbl = 4092;
    1752: ytbl = 4092;
    1753: ytbl = 4092;
    1754: ytbl = 4092;
    1755: ytbl = 4092;
    1756: ytbl = 4092;
    1757: ytbl = 4092;
    1758: ytbl = 4092;
    1759: ytbl = 4092;
    1760: ytbl = 4092;
    1761: ytbl = 4092;
    1762: ytbl = 4092;
    1763: ytbl = 4092;
    1764: ytbl = 4092;
    1765: ytbl = 4092;
    1766: ytbl = 4092;
    1767: ytbl = 4092;
    1768: ytbl = 4092;
    1769: ytbl = 4092;
    1770: ytbl = 4092;
    1771: ytbl = 4092;
    1772: ytbl = 4092;
    1773: ytbl = 4092;
    1774: ytbl = 4092;
    1775: ytbl = 4092;
    1776: ytbl = 4092;
    1777: ytbl = 4092;
    1778: ytbl = 4092;
    1779: ytbl = 4092;
    1780: ytbl = 4092;
    1781: ytbl = 4092;
    1782: ytbl = 4092;
    1783: ytbl = 4092;
    1784: ytbl = 4092;
    1785: ytbl = 4092;
    1786: ytbl = 4092;
    1787: ytbl = 4092;
    1788: ytbl = 4092;
    1789: ytbl = 4092;
    1790: ytbl = 4092;
    1791: ytbl = 4092;
    1792: ytbl = 4092;
    1793: ytbl = 4092;
    1794: ytbl = 4092;
    1795: ytbl = 4092;
    1796: ytbl = 4092;
    1797: ytbl = 4092;
    1798: ytbl = 4092;
    1799: ytbl = 4092;
    1800: ytbl = 4092;
    1801: ytbl = 4092;
    1802: ytbl = 4092;
    1803: ytbl = 4092;
    1804: ytbl = 4092;
    1805: ytbl = 4092;
    1806: ytbl = 4092;
    1807: ytbl = 4092;
    1808: ytbl = 4092;
    1809: ytbl = 4093;
    1810: ytbl = 4093;
    1811: ytbl = 4093;
    1812: ytbl = 4093;
    1813: ytbl = 4093;
    1814: ytbl = 4093;
    1815: ytbl = 4093;
    1816: ytbl = 4093;
    1817: ytbl = 4093;
    1818: ytbl = 4093;
    1819: ytbl = 4093;
    1820: ytbl = 4093;
    1821: ytbl = 4093;
    1822: ytbl = 4093;
    1823: ytbl = 4093;
    1824: ytbl = 4093;
    1825: ytbl = 4093;
    1826: ytbl = 4093;
    1827: ytbl = 4093;
    1828: ytbl = 4093;
    1829: ytbl = 4093;
    1830: ytbl = 4093;
    1831: ytbl = 4093;
    1832: ytbl = 4093;
    1833: ytbl = 4093;
    1834: ytbl = 4093;
    1835: ytbl = 4093;
    1836: ytbl = 4093;
    1837: ytbl = 4093;
    1838: ytbl = 4093;
    1839: ytbl = 4093;
    1840: ytbl = 4093;
    1841: ytbl = 4093;
    1842: ytbl = 4093;
    1843: ytbl = 4093;
    1844: ytbl = 4093;
    1845: ytbl = 4093;
    1846: ytbl = 4093;
    1847: ytbl = 4093;
    1848: ytbl = 4093;
    1849: ytbl = 4093;
    1850: ytbl = 4093;
    1851: ytbl = 4093;
    1852: ytbl = 4093;
    1853: ytbl = 4093;
    1854: ytbl = 4093;
    1855: ytbl = 4093;
    1856: ytbl = 4093;
    1857: ytbl = 4093;
    1858: ytbl = 4093;
    1859: ytbl = 4093;
    1860: ytbl = 4093;
    1861: ytbl = 4093;
    1862: ytbl = 4093;
    1863: ytbl = 4093;
    1864: ytbl = 4093;
    1865: ytbl = 4093;
    1866: ytbl = 4093;
    1867: ytbl = 4093;
    1868: ytbl = 4093;
    1869: ytbl = 4093;
    1870: ytbl = 4093;
    1871: ytbl = 4093;
    1872: ytbl = 4093;
    1873: ytbl = 4093;
    1874: ytbl = 4093;
    1875: ytbl = 4093;
    1876: ytbl = 4093;
    1877: ytbl = 4093;
    1878: ytbl = 4093;
    1879: ytbl = 4093;
    1880: ytbl = 4093;
    1881: ytbl = 4093;
    1882: ytbl = 4093;
    1883: ytbl = 4093;
    1884: ytbl = 4093;
    1885: ytbl = 4093;
    1886: ytbl = 4093;
    1887: ytbl = 4093;
    1888: ytbl = 4093;
    1889: ytbl = 4093;
    1890: ytbl = 4093;
    1891: ytbl = 4093;
    1892: ytbl = 4093;
    1893: ytbl = 4093;
    1894: ytbl = 4093;
    1895: ytbl = 4094;
    1896: ytbl = 4094;
    1897: ytbl = 4094;
    1898: ytbl = 4094;
    1899: ytbl = 4094;
    1900: ytbl = 4094;
    1901: ytbl = 4094;
    1902: ytbl = 4094;
    1903: ytbl = 4094;
    1904: ytbl = 4094;
    1905: ytbl = 4094;
    1906: ytbl = 4094;
    1907: ytbl = 4094;
    1908: ytbl = 4094;
    1909: ytbl = 4094;
    1910: ytbl = 4094;
    1911: ytbl = 4094;
    1912: ytbl = 4094;
    1913: ytbl = 4094;
    1914: ytbl = 4094;
    1915: ytbl = 4094;
    1916: ytbl = 4094;
    1917: ytbl = 4094;
    1918: ytbl = 4094;
    1919: ytbl = 4094;
    1920: ytbl = 4094;
    1921: ytbl = 4094;
    1922: ytbl = 4094;
    1923: ytbl = 4094;
    1924: ytbl = 4094;
    1925: ytbl = 4094;
    1926: ytbl = 4094;
    1927: ytbl = 4094;
    1928: ytbl = 4094;
    1929: ytbl = 4094;
    1930: ytbl = 4094;
    1931: ytbl = 4094;
    1932: ytbl = 4094;
    1933: ytbl = 4094;
    1934: ytbl = 4094;
    1935: ytbl = 4094;
    1936: ytbl = 4094;
    1937: ytbl = 4094;
    1938: ytbl = 4094;
    1939: ytbl = 4094;
    1940: ytbl = 4094;
    1941: ytbl = 4094;
    1942: ytbl = 4094;
    1943: ytbl = 4094;
    1944: ytbl = 4094;
    1945: ytbl = 4094;
    1946: ytbl = 4094;
    1947: ytbl = 4094;
    1948: ytbl = 4094;
    1949: ytbl = 4094;
    1950: ytbl = 4094;
    1951: ytbl = 4094;
    1952: ytbl = 4094;
    1953: ytbl = 4094;
    1954: ytbl = 4094;
    1955: ytbl = 4094;
    1956: ytbl = 4094;
    1957: ytbl = 4094;
    1958: ytbl = 4094;
    1959: ytbl = 4094;
    1960: ytbl = 4094;
    1961: ytbl = 4094;
    1962: ytbl = 4094;
    1963: ytbl = 4094;
    1964: ytbl = 4094;
    1965: ytbl = 4094;
    1966: ytbl = 4094;
    1967: ytbl = 4094;
    1968: ytbl = 4094;
    1969: ytbl = 4094;
    1970: ytbl = 4094;
    1971: ytbl = 4094;
    1972: ytbl = 4094;
    1973: ytbl = 4094;
    1974: ytbl = 4094;
    1975: ytbl = 4094;
    1976: ytbl = 4094;
    1977: ytbl = 4094;
    1978: ytbl = 4094;
    1979: ytbl = 4094;
    1980: ytbl = 4094;
    1981: ytbl = 4094;
    1982: ytbl = 4094;
    1983: ytbl = 4094;
    1984: ytbl = 4094;
    1985: ytbl = 4094;
    1986: ytbl = 4094;
    1987: ytbl = 4094;
    1988: ytbl = 4094;
    1989: ytbl = 4094;
    1990: ytbl = 4094;
    1991: ytbl = 4094;
    1992: ytbl = 4094;
    1993: ytbl = 4094;
    1994: ytbl = 4094;
    1995: ytbl = 4094;
    1996: ytbl = 4094;
    1997: ytbl = 4094;
    1998: ytbl = 4094;
    1999: ytbl = 4094;
    2000: ytbl = 4094;
    2001: ytbl = 4094;
    2002: ytbl = 4094;
    2003: ytbl = 4094;
    2004: ytbl = 4094;
    2005: ytbl = 4094;
    2006: ytbl = 4094;
    2007: ytbl = 4094;
    2008: ytbl = 4094;
    2009: ytbl = 4094;
    2010: ytbl = 4094;
    2011: ytbl = 4094;
    2012: ytbl = 4094;
    2013: ytbl = 4094;
    2014: ytbl = 4094;
    2015: ytbl = 4094;
    2016: ytbl = 4094;
    2017: ytbl = 4094;
    2018: ytbl = 4094;
    2019: ytbl = 4094;
    2020: ytbl = 4094;
    2021: ytbl = 4094;
    2022: ytbl = 4094;
    2023: ytbl = 4094;
    2024: ytbl = 4094;
    2025: ytbl = 4094;
    2026: ytbl = 4095;
    2027: ytbl = 4095;
    2028: ytbl = 4095;
    2029: ytbl = 4095;
    2030: ytbl = 4095;
    2031: ytbl = 4095;
    2032: ytbl = 4095;
    2033: ytbl = 4095;
    2034: ytbl = 4095;
    2035: ytbl = 4095;
    2036: ytbl = 4095;
    2037: ytbl = 4095;
    2038: ytbl = 4095;
    2039: ytbl = 4095;
    2040: ytbl = 4095;
    2041: ytbl = 4095;
    2042: ytbl = 4095;
    2043: ytbl = 4095;
    2044: ytbl = 4095;
    2045: ytbl = 4095;
    2046: ytbl = 4095;
    2047: ytbl = 4095;
    default: ytbl = 4095;
    endcase
end
endmodule
